VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 478.945 BY 489.665 ;
  PIN DataAdr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END DataAdr[0]
  PIN DataAdr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 485.665 228.990 489.665 ;
    END
  END DataAdr[10]
  PIN DataAdr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 469.240 478.945 469.840 ;
    END
  END DataAdr[11]
  PIN DataAdr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.808200 ;
    ANTENNADIFFAREA 1.918700 ;
    PORT
      LAYER met3 ;
        RECT 474.945 397.840 478.945 398.440 ;
    END
  END DataAdr[12]
  PIN DataAdr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 485.665 277.290 489.665 ;
    END
  END DataAdr[13]
  PIN DataAdr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END DataAdr[14]
  PIN DataAdr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met2 ;
        RECT 425.130 485.665 425.410 489.665 ;
    END
  END DataAdr[15]
  PIN DataAdr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 1.484000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END DataAdr[16]
  PIN DataAdr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER met3 ;
        RECT 474.945 17.040 478.945 17.640 ;
    END
  END DataAdr[17]
  PIN DataAdr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    ANTENNADIFFAREA 1.484000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 485.665 286.950 489.665 ;
    END
  END DataAdr[18]
  PIN DataAdr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 139.440 478.945 140.040 ;
    END
  END DataAdr[19]
  PIN DataAdr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 275.440 478.945 276.040 ;
    END
  END DataAdr[1]
  PIN DataAdr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 485.665 161.370 489.665 ;
    END
  END DataAdr[20]
  PIN DataAdr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END DataAdr[21]
  PIN DataAdr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER met2 ;
        RECT 206.170 485.665 206.450 489.665 ;
    END
  END DataAdr[22]
  PIN DataAdr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 1.484000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END DataAdr[23]
  PIN DataAdr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.342400 ;
    ANTENNADIFFAREA 8.078400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END DataAdr[24]
  PIN DataAdr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END DataAdr[25]
  PIN DataAdr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER met3 ;
        RECT 474.945 224.440 478.945 225.040 ;
    END
  END DataAdr[26]
  PIN DataAdr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 485.665 45.450 489.665 ;
    END
  END DataAdr[27]
  PIN DataAdr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 485.665 322.370 489.665 ;
    END
  END DataAdr[28]
  PIN DataAdr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END DataAdr[29]
  PIN DataAdr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END DataAdr[2]
  PIN DataAdr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met2 ;
        RECT 473.430 485.665 473.710 489.665 ;
    END
  END DataAdr[30]
  PIN DataAdr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END DataAdr[31]
  PIN DataAdr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END DataAdr[3]
  PIN DataAdr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 54.440 478.945 55.040 ;
    END
  END DataAdr[4]
  PIN DataAdr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.603600 ;
    ANTENNADIFFAREA 4.814100 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END DataAdr[5]
  PIN DataAdr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 2.090400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END DataAdr[6]
  PIN DataAdr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END DataAdr[7]
  PIN DataAdr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END DataAdr[8]
  PIN DataAdr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 1.484000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 485.665 125.950 489.665 ;
    END
  END DataAdr[9]
  PIN Instr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.848500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 485.665 264.410 489.665 ;
    END
  END Instr[0]
  PIN Instr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.081500 ;
    PORT
      LAYER met2 ;
        RECT 438.010 485.665 438.290 489.665 ;
    END
  END Instr[10]
  PIN Instr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.198400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END Instr[11]
  PIN Instr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 485.665 55.110 489.665 ;
    END
  END Instr[12]
  PIN Instr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.494000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 384.240 478.945 384.840 ;
    END
  END Instr[13]
  PIN Instr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.363500 ;
    PORT
      LAYER met2 ;
        RECT 460.550 485.665 460.830 489.665 ;
    END
  END Instr[14]
  PIN Instr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.663500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 360.440 478.945 361.040 ;
    END
  END Instr[15]
  PIN Instr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611900 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END Instr[16]
  PIN Instr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.830000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END Instr[17]
  PIN Instr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END Instr[18]
  PIN Instr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.469500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 200.640 478.945 201.240 ;
    END
  END Instr[19]
  PIN Instr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.848500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END Instr[1]
  PIN Instr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.089500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END Instr[20]
  PIN Instr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.597300 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 474.945 30.640 478.945 31.240 ;
    END
  END Instr[21]
  PIN Instr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.047000 ;
    PORT
      LAYER met2 ;
        RECT 183.630 485.665 183.910 489.665 ;
    END
  END Instr[22]
  PIN Instr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END Instr[23]
  PIN Instr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END Instr[24]
  PIN Instr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.601000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END Instr[25]
  PIN Instr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 485.665 219.330 489.665 ;
    END
  END Instr[26]
  PIN Instr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 485.665 32.570 489.665 ;
    END
  END Instr[27]
  PIN Instr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.611000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 370.640 478.945 371.240 ;
    END
  END Instr[28]
  PIN Instr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.177100 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END Instr[29]
  PIN Instr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.197500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END Instr[2]
  PIN Instr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.984500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 485.665 171.030 489.665 ;
    END
  END Instr[30]
  PIN Instr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.823500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 115.640 478.945 116.240 ;
    END
  END Instr[31]
  PIN Instr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.197500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 421.640 478.945 422.240 ;
    END
  END Instr[3]
  PIN Instr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.950000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 163.240 478.945 163.840 ;
    END
  END Instr[4]
  PIN Instr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.465000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END Instr[5]
  PIN Instr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 64.640 478.945 65.240 ;
    END
  END Instr[6]
  PIN Instr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.449500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END Instr[7]
  PIN Instr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.532800 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END Instr[8]
  PIN Instr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.208400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 474.945 445.440 478.945 446.040 ;
    END
  END Instr[9]
  PIN MemWrite
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END MemWrite
  PIN PC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.560000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 450.890 485.665 451.170 489.665 ;
    END
  END PC[0]
  PIN PC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.853000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END PC[10]
  PIN PC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.368000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END PC[11]
  PIN PC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.863000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 334.970 485.665 335.250 489.665 ;
    END
  END PC[12]
  PIN PC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 309.210 485.665 309.490 489.665 ;
    END
  END PC[13]
  PIN PC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.731500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 485.665 148.490 489.665 ;
    END
  END PC[14]
  PIN PC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END PC[15]
  PIN PC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 485.665 19.690 489.665 ;
    END
  END PC[16]
  PIN PC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 431.840 478.945 432.440 ;
    END
  END PC[17]
  PIN PC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.737000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END PC[18]
  PIN PC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.489500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END PC[19]
  PIN PC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 346.840 478.945 347.440 ;
    END
  END PC[1]
  PIN PC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.620000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END PC[20]
  PIN PC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.863000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END PC[21]
  PIN PC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.120500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 299.240 478.945 299.840 ;
    END
  END PC[22]
  PIN PC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.853000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END PC[23]
  PIN PC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 102.040 478.945 102.640 ;
    END
  END PC[24]
  PIN PC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.727000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 485.665 113.070 489.665 ;
    END
  END PC[25]
  PIN PC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.615500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 187.040 478.945 187.640 ;
    END
  END PC[26]
  PIN PC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.242000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END PC[27]
  PIN PC[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.727000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 415.470 485.665 415.750 489.665 ;
    END
  END PC[28]
  PIN PC[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.601000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 214.240 478.945 214.840 ;
    END
  END PC[29]
  PIN PC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.339000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END PC[2]
  PIN PC[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.984500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END PC[30]
  PIN PC[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.242000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 485.665 299.830 489.665 ;
    END
  END PC[31]
  PIN PC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.343500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END PC[3]
  PIN PC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.858500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END PC[4]
  PIN PC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.285000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 485.665 10.030 489.665 ;
    END
  END PC[5]
  PIN PC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.368000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 485.665 67.990 489.665 ;
    END
  END PC[6]
  PIN PC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.994500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 367.170 485.665 367.450 489.665 ;
    END
  END PC[7]
  PIN PC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.232000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 485.665 380.330 489.665 ;
    END
  END PC[8]
  PIN PC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.873000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 485.665 357.790 489.665 ;
    END
  END PC[9]
  PIN ReadData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.907700 ;
    ANTENNADIFFAREA 4.781700 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END ReadData[0]
  PIN ReadData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END ReadData[10]
  PIN ReadData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 474.945 40.840 478.945 41.440 ;
    END
  END ReadData[11]
  PIN ReadData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.299500 ;
    ANTENNADIFFAREA 2.173500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END ReadData[12]
  PIN ReadData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.330 485.665 135.610 489.665 ;
    END
  END ReadData[13]
  PIN ReadData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 248.240 478.945 248.840 ;
    END
  END ReadData[14]
  PIN ReadData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 392.930 485.665 393.210 489.665 ;
    END
  END ReadData[15]
  PIN ReadData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END ReadData[16]
  PIN ReadData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.168900 ;
    ANTENNADIFFAREA 3.042900 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END ReadData[17]
  PIN ReadData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 261.840 478.945 262.440 ;
    END
  END ReadData[18]
  PIN ReadData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 193.290 485.665 193.570 489.665 ;
    END
  END ReadData[19]
  PIN ReadData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 176.840 478.945 177.440 ;
    END
  END ReadData[1]
  PIN ReadData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END ReadData[20]
  PIN ReadData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.116900 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END ReadData[21]
  PIN ReadData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 336.640 478.945 337.240 ;
    END
  END ReadData[22]
  PIN ReadData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END ReadData[23]
  PIN ReadData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.603600 ;
    ANTENNADIFFAREA 3.477600 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END ReadData[24]
  PIN ReadData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 474.945 125.840 478.945 126.440 ;
    END
  END ReadData[25]
  PIN ReadData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END ReadData[26]
  PIN ReadData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 474.945 3.440 478.945 4.040 ;
    END
  END ReadData[27]
  PIN ReadData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 103.130 485.665 103.410 489.665 ;
    END
  END ReadData[28]
  PIN ReadData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END ReadData[29]
  PIN ReadData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END ReadData[2]
  PIN ReadData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END ReadData[30]
  PIN ReadData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 474.945 78.240 478.945 78.840 ;
    END
  END ReadData[31]
  PIN ReadData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 474.945 408.040 478.945 408.640 ;
    END
  END ReadData[3]
  PIN ReadData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 285.640 478.945 286.240 ;
    END
  END ReadData[4]
  PIN ReadData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.473000 ;
    ANTENNADIFFAREA 4.347000 ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END ReadData[5]
  PIN ReadData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END ReadData[6]
  PIN ReadData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 474.945 153.040 478.945 153.640 ;
    END
  END ReadData[7]
  PIN ReadData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END ReadData[8]
  PIN ReadData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 309.440 478.945 310.040 ;
    END
  END ReadData[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 478.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 478.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 478.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 473.580 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 473.580 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 473.580 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 478.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 478.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 478.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 473.580 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 473.580 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 473.580 334.690 ;
    END
  END VPWR
  PIN WriteData[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 474.945 459.040 478.945 459.640 ;
    END
  END WriteData[0]
  PIN WriteData[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END WriteData[10]
  PIN WriteData[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 482.840 478.945 483.440 ;
    END
  END WriteData[11]
  PIN WriteData[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END WriteData[12]
  PIN WriteData[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END WriteData[13]
  PIN WriteData[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END WriteData[14]
  PIN WriteData[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END WriteData[15]
  PIN WriteData[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END WriteData[16]
  PIN WriteData[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END WriteData[17]
  PIN WriteData[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 485.665 90.530 489.665 ;
    END
  END WriteData[18]
  PIN WriteData[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 485.665 251.530 489.665 ;
    END
  END WriteData[19]
  PIN WriteData[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END WriteData[1]
  PIN WriteData[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END WriteData[20]
  PIN WriteData[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END WriteData[21]
  PIN WriteData[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END WriteData[22]
  PIN WriteData[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 241.590 485.665 241.870 489.665 ;
    END
  END WriteData[23]
  PIN WriteData[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END WriteData[24]
  PIN WriteData[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.911000 ;
    PORT
      LAYER met2 ;
        RECT 402.590 485.665 402.870 489.665 ;
    END
  END WriteData[25]
  PIN WriteData[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 91.840 478.945 92.440 ;
    END
  END WriteData[26]
  PIN WriteData[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END WriteData[27]
  PIN WriteData[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END WriteData[28]
  PIN WriteData[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.911000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END WriteData[29]
  PIN WriteData[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END WriteData[2]
  PIN WriteData[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.911000 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END WriteData[30]
  PIN WriteData[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 474.945 323.040 478.945 323.640 ;
    END
  END WriteData[31]
  PIN WriteData[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END WriteData[3]
  PIN WriteData[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END WriteData[4]
  PIN WriteData[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 344.630 485.665 344.910 489.665 ;
    END
  END WriteData[5]
  PIN WriteData[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END WriteData[6]
  PIN WriteData[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 485.665 77.650 489.665 ;
    END
  END WriteData[7]
  PIN WriteData[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END WriteData[8]
  PIN WriteData[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END WriteData[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.732500 ;
    PORT
      LAYER met3 ;
        RECT 474.945 238.040 478.945 238.640 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 473.340 478.805 ;
      LAYER met1 ;
        RECT 4.670 10.640 473.730 478.960 ;
      LAYER met2 ;
        RECT 0.090 485.385 9.470 486.725 ;
        RECT 10.310 485.385 19.130 486.725 ;
        RECT 19.970 485.385 32.010 486.725 ;
        RECT 32.850 485.385 44.890 486.725 ;
        RECT 45.730 485.385 54.550 486.725 ;
        RECT 55.390 485.385 67.430 486.725 ;
        RECT 68.270 485.385 77.090 486.725 ;
        RECT 77.930 485.385 89.970 486.725 ;
        RECT 90.810 485.385 102.850 486.725 ;
        RECT 103.690 485.385 112.510 486.725 ;
        RECT 113.350 485.385 125.390 486.725 ;
        RECT 126.230 485.385 135.050 486.725 ;
        RECT 135.890 485.385 147.930 486.725 ;
        RECT 148.770 485.385 160.810 486.725 ;
        RECT 161.650 485.385 170.470 486.725 ;
        RECT 171.310 485.385 183.350 486.725 ;
        RECT 184.190 485.385 193.010 486.725 ;
        RECT 193.850 485.385 205.890 486.725 ;
        RECT 206.730 485.385 218.770 486.725 ;
        RECT 219.610 485.385 228.430 486.725 ;
        RECT 229.270 485.385 241.310 486.725 ;
        RECT 242.150 485.385 250.970 486.725 ;
        RECT 251.810 485.385 263.850 486.725 ;
        RECT 264.690 485.385 276.730 486.725 ;
        RECT 277.570 485.385 286.390 486.725 ;
        RECT 287.230 485.385 299.270 486.725 ;
        RECT 300.110 485.385 308.930 486.725 ;
        RECT 309.770 485.385 321.810 486.725 ;
        RECT 322.650 485.385 334.690 486.725 ;
        RECT 335.530 485.385 344.350 486.725 ;
        RECT 345.190 485.385 357.230 486.725 ;
        RECT 358.070 485.385 366.890 486.725 ;
        RECT 367.730 485.385 379.770 486.725 ;
        RECT 380.610 485.385 392.650 486.725 ;
        RECT 393.490 485.385 402.310 486.725 ;
        RECT 403.150 485.385 415.190 486.725 ;
        RECT 416.030 485.385 424.850 486.725 ;
        RECT 425.690 485.385 437.730 486.725 ;
        RECT 438.570 485.385 450.610 486.725 ;
        RECT 451.450 485.385 460.270 486.725 ;
        RECT 461.110 485.385 473.150 486.725 ;
        RECT 0.090 4.280 473.710 485.385 ;
        RECT 0.650 3.670 9.470 4.280 ;
        RECT 10.310 3.670 22.350 4.280 ;
        RECT 23.190 3.670 32.010 4.280 ;
        RECT 32.850 3.670 44.890 4.280 ;
        RECT 45.730 3.670 54.550 4.280 ;
        RECT 55.390 3.670 67.430 4.280 ;
        RECT 68.270 3.670 80.310 4.280 ;
        RECT 81.150 3.670 89.970 4.280 ;
        RECT 90.810 3.670 102.850 4.280 ;
        RECT 103.690 3.670 112.510 4.280 ;
        RECT 113.350 3.670 125.390 4.280 ;
        RECT 126.230 3.670 138.270 4.280 ;
        RECT 139.110 3.670 147.930 4.280 ;
        RECT 148.770 3.670 160.810 4.280 ;
        RECT 161.650 3.670 170.470 4.280 ;
        RECT 171.310 3.670 183.350 4.280 ;
        RECT 184.190 3.670 196.230 4.280 ;
        RECT 197.070 3.670 205.890 4.280 ;
        RECT 206.730 3.670 218.770 4.280 ;
        RECT 219.610 3.670 228.430 4.280 ;
        RECT 229.270 3.670 241.310 4.280 ;
        RECT 242.150 3.670 254.190 4.280 ;
        RECT 255.030 3.670 263.850 4.280 ;
        RECT 264.690 3.670 276.730 4.280 ;
        RECT 277.570 3.670 286.390 4.280 ;
        RECT 287.230 3.670 299.270 4.280 ;
        RECT 300.110 3.670 312.150 4.280 ;
        RECT 312.990 3.670 321.810 4.280 ;
        RECT 322.650 3.670 334.690 4.280 ;
        RECT 335.530 3.670 344.350 4.280 ;
        RECT 345.190 3.670 357.230 4.280 ;
        RECT 358.070 3.670 370.110 4.280 ;
        RECT 370.950 3.670 379.770 4.280 ;
        RECT 380.610 3.670 392.650 4.280 ;
        RECT 393.490 3.670 402.310 4.280 ;
        RECT 403.150 3.670 415.190 4.280 ;
        RECT 416.030 3.670 428.070 4.280 ;
        RECT 428.910 3.670 437.730 4.280 ;
        RECT 438.570 3.670 450.610 4.280 ;
        RECT 451.450 3.670 460.270 4.280 ;
        RECT 461.110 3.670 473.150 4.280 ;
      LAYER met3 ;
        RECT 4.400 485.840 475.330 486.705 ;
        RECT 0.065 483.840 475.330 485.840 ;
        RECT 0.065 482.440 474.545 483.840 ;
        RECT 0.065 477.040 475.330 482.440 ;
        RECT 4.400 475.640 475.330 477.040 ;
        RECT 0.065 470.240 475.330 475.640 ;
        RECT 0.065 468.840 474.545 470.240 ;
        RECT 0.065 463.440 475.330 468.840 ;
        RECT 4.400 462.040 475.330 463.440 ;
        RECT 0.065 460.040 475.330 462.040 ;
        RECT 0.065 458.640 474.545 460.040 ;
        RECT 0.065 453.240 475.330 458.640 ;
        RECT 4.400 451.840 475.330 453.240 ;
        RECT 0.065 446.440 475.330 451.840 ;
        RECT 0.065 445.040 474.545 446.440 ;
        RECT 0.065 439.640 475.330 445.040 ;
        RECT 4.400 438.240 475.330 439.640 ;
        RECT 0.065 432.840 475.330 438.240 ;
        RECT 0.065 431.440 474.545 432.840 ;
        RECT 0.065 426.040 475.330 431.440 ;
        RECT 4.400 424.640 475.330 426.040 ;
        RECT 0.065 422.640 475.330 424.640 ;
        RECT 0.065 421.240 474.545 422.640 ;
        RECT 0.065 415.840 475.330 421.240 ;
        RECT 4.400 414.440 475.330 415.840 ;
        RECT 0.065 409.040 475.330 414.440 ;
        RECT 0.065 407.640 474.545 409.040 ;
        RECT 0.065 402.240 475.330 407.640 ;
        RECT 4.400 400.840 475.330 402.240 ;
        RECT 0.065 398.840 475.330 400.840 ;
        RECT 0.065 397.440 474.545 398.840 ;
        RECT 0.065 392.040 475.330 397.440 ;
        RECT 4.400 390.640 475.330 392.040 ;
        RECT 0.065 385.240 475.330 390.640 ;
        RECT 0.065 383.840 474.545 385.240 ;
        RECT 0.065 378.440 475.330 383.840 ;
        RECT 4.400 377.040 475.330 378.440 ;
        RECT 0.065 371.640 475.330 377.040 ;
        RECT 0.065 370.240 474.545 371.640 ;
        RECT 0.065 364.840 475.330 370.240 ;
        RECT 4.400 363.440 475.330 364.840 ;
        RECT 0.065 361.440 475.330 363.440 ;
        RECT 0.065 360.040 474.545 361.440 ;
        RECT 0.065 354.640 475.330 360.040 ;
        RECT 4.400 353.240 475.330 354.640 ;
        RECT 0.065 347.840 475.330 353.240 ;
        RECT 0.065 346.440 474.545 347.840 ;
        RECT 0.065 341.040 475.330 346.440 ;
        RECT 4.400 339.640 475.330 341.040 ;
        RECT 0.065 337.640 475.330 339.640 ;
        RECT 0.065 336.240 474.545 337.640 ;
        RECT 0.065 330.840 475.330 336.240 ;
        RECT 4.400 329.440 475.330 330.840 ;
        RECT 0.065 324.040 475.330 329.440 ;
        RECT 0.065 322.640 474.545 324.040 ;
        RECT 0.065 317.240 475.330 322.640 ;
        RECT 4.400 315.840 475.330 317.240 ;
        RECT 0.065 310.440 475.330 315.840 ;
        RECT 0.065 309.040 474.545 310.440 ;
        RECT 0.065 303.640 475.330 309.040 ;
        RECT 4.400 302.240 475.330 303.640 ;
        RECT 0.065 300.240 475.330 302.240 ;
        RECT 0.065 298.840 474.545 300.240 ;
        RECT 0.065 293.440 475.330 298.840 ;
        RECT 4.400 292.040 475.330 293.440 ;
        RECT 0.065 286.640 475.330 292.040 ;
        RECT 0.065 285.240 474.545 286.640 ;
        RECT 0.065 279.840 475.330 285.240 ;
        RECT 4.400 278.440 475.330 279.840 ;
        RECT 0.065 276.440 475.330 278.440 ;
        RECT 0.065 275.040 474.545 276.440 ;
        RECT 0.065 269.640 475.330 275.040 ;
        RECT 4.400 268.240 475.330 269.640 ;
        RECT 0.065 262.840 475.330 268.240 ;
        RECT 0.065 261.440 474.545 262.840 ;
        RECT 0.065 256.040 475.330 261.440 ;
        RECT 4.400 254.640 475.330 256.040 ;
        RECT 0.065 249.240 475.330 254.640 ;
        RECT 0.065 247.840 474.545 249.240 ;
        RECT 0.065 242.440 475.330 247.840 ;
        RECT 4.400 241.040 475.330 242.440 ;
        RECT 0.065 239.040 475.330 241.040 ;
        RECT 0.065 237.640 474.545 239.040 ;
        RECT 0.065 232.240 475.330 237.640 ;
        RECT 4.400 230.840 475.330 232.240 ;
        RECT 0.065 225.440 475.330 230.840 ;
        RECT 0.065 224.040 474.545 225.440 ;
        RECT 0.065 218.640 475.330 224.040 ;
        RECT 4.400 217.240 475.330 218.640 ;
        RECT 0.065 215.240 475.330 217.240 ;
        RECT 0.065 213.840 474.545 215.240 ;
        RECT 0.065 208.440 475.330 213.840 ;
        RECT 4.400 207.040 475.330 208.440 ;
        RECT 0.065 201.640 475.330 207.040 ;
        RECT 0.065 200.240 474.545 201.640 ;
        RECT 0.065 194.840 475.330 200.240 ;
        RECT 4.400 193.440 475.330 194.840 ;
        RECT 0.065 188.040 475.330 193.440 ;
        RECT 0.065 186.640 474.545 188.040 ;
        RECT 0.065 181.240 475.330 186.640 ;
        RECT 4.400 179.840 475.330 181.240 ;
        RECT 0.065 177.840 475.330 179.840 ;
        RECT 0.065 176.440 474.545 177.840 ;
        RECT 0.065 171.040 475.330 176.440 ;
        RECT 4.400 169.640 475.330 171.040 ;
        RECT 0.065 164.240 475.330 169.640 ;
        RECT 0.065 162.840 474.545 164.240 ;
        RECT 0.065 157.440 475.330 162.840 ;
        RECT 4.400 156.040 475.330 157.440 ;
        RECT 0.065 154.040 475.330 156.040 ;
        RECT 0.065 152.640 474.545 154.040 ;
        RECT 0.065 147.240 475.330 152.640 ;
        RECT 4.400 145.840 475.330 147.240 ;
        RECT 0.065 140.440 475.330 145.840 ;
        RECT 0.065 139.040 474.545 140.440 ;
        RECT 0.065 133.640 475.330 139.040 ;
        RECT 4.400 132.240 475.330 133.640 ;
        RECT 0.065 126.840 475.330 132.240 ;
        RECT 0.065 125.440 474.545 126.840 ;
        RECT 0.065 120.040 475.330 125.440 ;
        RECT 4.400 118.640 475.330 120.040 ;
        RECT 0.065 116.640 475.330 118.640 ;
        RECT 0.065 115.240 474.545 116.640 ;
        RECT 0.065 109.840 475.330 115.240 ;
        RECT 4.400 108.440 475.330 109.840 ;
        RECT 0.065 103.040 475.330 108.440 ;
        RECT 0.065 101.640 474.545 103.040 ;
        RECT 0.065 96.240 475.330 101.640 ;
        RECT 4.400 94.840 475.330 96.240 ;
        RECT 0.065 92.840 475.330 94.840 ;
        RECT 0.065 91.440 474.545 92.840 ;
        RECT 0.065 86.040 475.330 91.440 ;
        RECT 4.400 84.640 475.330 86.040 ;
        RECT 0.065 79.240 475.330 84.640 ;
        RECT 0.065 77.840 474.545 79.240 ;
        RECT 0.065 72.440 475.330 77.840 ;
        RECT 4.400 71.040 475.330 72.440 ;
        RECT 0.065 65.640 475.330 71.040 ;
        RECT 0.065 64.240 474.545 65.640 ;
        RECT 0.065 58.840 475.330 64.240 ;
        RECT 4.400 57.440 475.330 58.840 ;
        RECT 0.065 55.440 475.330 57.440 ;
        RECT 0.065 54.040 474.545 55.440 ;
        RECT 0.065 48.640 475.330 54.040 ;
        RECT 4.400 47.240 475.330 48.640 ;
        RECT 0.065 41.840 475.330 47.240 ;
        RECT 0.065 40.440 474.545 41.840 ;
        RECT 0.065 35.040 475.330 40.440 ;
        RECT 4.400 33.640 475.330 35.040 ;
        RECT 0.065 31.640 475.330 33.640 ;
        RECT 0.065 30.240 474.545 31.640 ;
        RECT 0.065 24.840 475.330 30.240 ;
        RECT 4.400 23.440 475.330 24.840 ;
        RECT 0.065 18.040 475.330 23.440 ;
        RECT 0.065 16.640 474.545 18.040 ;
        RECT 0.065 11.240 475.330 16.640 ;
        RECT 4.400 9.840 475.330 11.240 ;
        RECT 0.065 4.440 475.330 9.840 ;
        RECT 0.065 3.580 474.545 4.440 ;
      LAYER met4 ;
        RECT 16.855 10.240 20.640 472.425 ;
        RECT 23.040 10.240 23.940 472.425 ;
        RECT 26.340 10.240 174.240 472.425 ;
        RECT 176.640 10.240 177.540 472.425 ;
        RECT 179.940 10.240 327.840 472.425 ;
        RECT 330.240 10.240 331.140 472.425 ;
        RECT 333.540 10.240 447.745 472.425 ;
        RECT 16.855 3.575 447.745 10.240 ;
  END
END top
END LIBRARY

