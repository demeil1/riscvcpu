module top (MemWrite,
    clk,
    reset,
    DataAdr,
    Instr,
    PC,
    ReadData,
    WriteData);
 output MemWrite;
 input clk;
 input reset;
 output [31:0] DataAdr;
 input [31:0] Instr;
 output [31:0] PC;
 input [31:0] ReadData;
 output [31:0] WriteData;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire \rvsingle.dp.PCNext[10] ;
 wire \rvsingle.dp.PCNext[11] ;
 wire \rvsingle.dp.PCNext[12] ;
 wire \rvsingle.dp.PCNext[13] ;
 wire \rvsingle.dp.PCNext[14] ;
 wire \rvsingle.dp.PCNext[15] ;
 wire \rvsingle.dp.PCNext[16] ;
 wire \rvsingle.dp.PCNext[17] ;
 wire \rvsingle.dp.PCNext[18] ;
 wire \rvsingle.dp.PCNext[19] ;
 wire \rvsingle.dp.PCNext[20] ;
 wire \rvsingle.dp.PCNext[21] ;
 wire \rvsingle.dp.PCNext[22] ;
 wire \rvsingle.dp.PCNext[23] ;
 wire \rvsingle.dp.PCNext[24] ;
 wire \rvsingle.dp.PCNext[25] ;
 wire \rvsingle.dp.PCNext[26] ;
 wire \rvsingle.dp.PCNext[27] ;
 wire \rvsingle.dp.PCNext[28] ;
 wire \rvsingle.dp.PCNext[29] ;
 wire \rvsingle.dp.PCNext[2] ;
 wire \rvsingle.dp.PCNext[30] ;
 wire \rvsingle.dp.PCNext[31] ;
 wire \rvsingle.dp.PCNext[3] ;
 wire \rvsingle.dp.PCNext[4] ;
 wire \rvsingle.dp.PCNext[5] ;
 wire \rvsingle.dp.PCNext[6] ;
 wire \rvsingle.dp.PCNext[7] ;
 wire \rvsingle.dp.PCNext[8] ;
 wire \rvsingle.dp.PCNext[9] ;
 wire \rvsingle.dp.rf.rf[0][0] ;
 wire \rvsingle.dp.rf.rf[0][10] ;
 wire \rvsingle.dp.rf.rf[0][11] ;
 wire \rvsingle.dp.rf.rf[0][12] ;
 wire \rvsingle.dp.rf.rf[0][13] ;
 wire \rvsingle.dp.rf.rf[0][14] ;
 wire \rvsingle.dp.rf.rf[0][15] ;
 wire \rvsingle.dp.rf.rf[0][16] ;
 wire \rvsingle.dp.rf.rf[0][17] ;
 wire \rvsingle.dp.rf.rf[0][18] ;
 wire \rvsingle.dp.rf.rf[0][19] ;
 wire \rvsingle.dp.rf.rf[0][1] ;
 wire \rvsingle.dp.rf.rf[0][20] ;
 wire \rvsingle.dp.rf.rf[0][21] ;
 wire \rvsingle.dp.rf.rf[0][22] ;
 wire \rvsingle.dp.rf.rf[0][23] ;
 wire \rvsingle.dp.rf.rf[0][24] ;
 wire \rvsingle.dp.rf.rf[0][25] ;
 wire \rvsingle.dp.rf.rf[0][26] ;
 wire \rvsingle.dp.rf.rf[0][27] ;
 wire \rvsingle.dp.rf.rf[0][28] ;
 wire \rvsingle.dp.rf.rf[0][29] ;
 wire \rvsingle.dp.rf.rf[0][2] ;
 wire \rvsingle.dp.rf.rf[0][30] ;
 wire \rvsingle.dp.rf.rf[0][31] ;
 wire \rvsingle.dp.rf.rf[0][3] ;
 wire \rvsingle.dp.rf.rf[0][4] ;
 wire \rvsingle.dp.rf.rf[0][5] ;
 wire \rvsingle.dp.rf.rf[0][6] ;
 wire \rvsingle.dp.rf.rf[0][7] ;
 wire \rvsingle.dp.rf.rf[0][8] ;
 wire \rvsingle.dp.rf.rf[0][9] ;
 wire \rvsingle.dp.rf.rf[10][0] ;
 wire \rvsingle.dp.rf.rf[10][10] ;
 wire \rvsingle.dp.rf.rf[10][11] ;
 wire \rvsingle.dp.rf.rf[10][12] ;
 wire \rvsingle.dp.rf.rf[10][13] ;
 wire \rvsingle.dp.rf.rf[10][14] ;
 wire \rvsingle.dp.rf.rf[10][15] ;
 wire \rvsingle.dp.rf.rf[10][16] ;
 wire \rvsingle.dp.rf.rf[10][17] ;
 wire \rvsingle.dp.rf.rf[10][18] ;
 wire \rvsingle.dp.rf.rf[10][19] ;
 wire \rvsingle.dp.rf.rf[10][1] ;
 wire \rvsingle.dp.rf.rf[10][20] ;
 wire \rvsingle.dp.rf.rf[10][21] ;
 wire \rvsingle.dp.rf.rf[10][22] ;
 wire \rvsingle.dp.rf.rf[10][23] ;
 wire \rvsingle.dp.rf.rf[10][24] ;
 wire \rvsingle.dp.rf.rf[10][25] ;
 wire \rvsingle.dp.rf.rf[10][26] ;
 wire \rvsingle.dp.rf.rf[10][27] ;
 wire \rvsingle.dp.rf.rf[10][28] ;
 wire \rvsingle.dp.rf.rf[10][29] ;
 wire \rvsingle.dp.rf.rf[10][2] ;
 wire \rvsingle.dp.rf.rf[10][30] ;
 wire \rvsingle.dp.rf.rf[10][31] ;
 wire \rvsingle.dp.rf.rf[10][3] ;
 wire \rvsingle.dp.rf.rf[10][4] ;
 wire \rvsingle.dp.rf.rf[10][5] ;
 wire \rvsingle.dp.rf.rf[10][6] ;
 wire \rvsingle.dp.rf.rf[10][7] ;
 wire \rvsingle.dp.rf.rf[10][8] ;
 wire \rvsingle.dp.rf.rf[10][9] ;
 wire \rvsingle.dp.rf.rf[11][0] ;
 wire \rvsingle.dp.rf.rf[11][10] ;
 wire \rvsingle.dp.rf.rf[11][11] ;
 wire \rvsingle.dp.rf.rf[11][12] ;
 wire \rvsingle.dp.rf.rf[11][13] ;
 wire \rvsingle.dp.rf.rf[11][14] ;
 wire \rvsingle.dp.rf.rf[11][15] ;
 wire \rvsingle.dp.rf.rf[11][16] ;
 wire \rvsingle.dp.rf.rf[11][17] ;
 wire \rvsingle.dp.rf.rf[11][18] ;
 wire \rvsingle.dp.rf.rf[11][19] ;
 wire \rvsingle.dp.rf.rf[11][1] ;
 wire \rvsingle.dp.rf.rf[11][20] ;
 wire \rvsingle.dp.rf.rf[11][21] ;
 wire \rvsingle.dp.rf.rf[11][22] ;
 wire \rvsingle.dp.rf.rf[11][23] ;
 wire \rvsingle.dp.rf.rf[11][24] ;
 wire \rvsingle.dp.rf.rf[11][25] ;
 wire \rvsingle.dp.rf.rf[11][26] ;
 wire \rvsingle.dp.rf.rf[11][27] ;
 wire \rvsingle.dp.rf.rf[11][28] ;
 wire \rvsingle.dp.rf.rf[11][29] ;
 wire \rvsingle.dp.rf.rf[11][2] ;
 wire \rvsingle.dp.rf.rf[11][30] ;
 wire \rvsingle.dp.rf.rf[11][31] ;
 wire \rvsingle.dp.rf.rf[11][3] ;
 wire \rvsingle.dp.rf.rf[11][4] ;
 wire \rvsingle.dp.rf.rf[11][5] ;
 wire \rvsingle.dp.rf.rf[11][6] ;
 wire \rvsingle.dp.rf.rf[11][7] ;
 wire \rvsingle.dp.rf.rf[11][8] ;
 wire \rvsingle.dp.rf.rf[11][9] ;
 wire \rvsingle.dp.rf.rf[12][0] ;
 wire \rvsingle.dp.rf.rf[12][10] ;
 wire \rvsingle.dp.rf.rf[12][11] ;
 wire \rvsingle.dp.rf.rf[12][12] ;
 wire \rvsingle.dp.rf.rf[12][13] ;
 wire \rvsingle.dp.rf.rf[12][14] ;
 wire \rvsingle.dp.rf.rf[12][15] ;
 wire \rvsingle.dp.rf.rf[12][16] ;
 wire \rvsingle.dp.rf.rf[12][17] ;
 wire \rvsingle.dp.rf.rf[12][18] ;
 wire \rvsingle.dp.rf.rf[12][19] ;
 wire \rvsingle.dp.rf.rf[12][1] ;
 wire \rvsingle.dp.rf.rf[12][20] ;
 wire \rvsingle.dp.rf.rf[12][21] ;
 wire \rvsingle.dp.rf.rf[12][22] ;
 wire \rvsingle.dp.rf.rf[12][23] ;
 wire \rvsingle.dp.rf.rf[12][24] ;
 wire \rvsingle.dp.rf.rf[12][25] ;
 wire \rvsingle.dp.rf.rf[12][26] ;
 wire \rvsingle.dp.rf.rf[12][27] ;
 wire \rvsingle.dp.rf.rf[12][28] ;
 wire \rvsingle.dp.rf.rf[12][29] ;
 wire \rvsingle.dp.rf.rf[12][2] ;
 wire \rvsingle.dp.rf.rf[12][30] ;
 wire \rvsingle.dp.rf.rf[12][31] ;
 wire \rvsingle.dp.rf.rf[12][3] ;
 wire \rvsingle.dp.rf.rf[12][4] ;
 wire \rvsingle.dp.rf.rf[12][5] ;
 wire \rvsingle.dp.rf.rf[12][6] ;
 wire \rvsingle.dp.rf.rf[12][7] ;
 wire \rvsingle.dp.rf.rf[12][8] ;
 wire \rvsingle.dp.rf.rf[12][9] ;
 wire \rvsingle.dp.rf.rf[13][0] ;
 wire \rvsingle.dp.rf.rf[13][10] ;
 wire \rvsingle.dp.rf.rf[13][11] ;
 wire \rvsingle.dp.rf.rf[13][12] ;
 wire \rvsingle.dp.rf.rf[13][13] ;
 wire \rvsingle.dp.rf.rf[13][14] ;
 wire \rvsingle.dp.rf.rf[13][15] ;
 wire \rvsingle.dp.rf.rf[13][16] ;
 wire \rvsingle.dp.rf.rf[13][17] ;
 wire \rvsingle.dp.rf.rf[13][18] ;
 wire \rvsingle.dp.rf.rf[13][19] ;
 wire \rvsingle.dp.rf.rf[13][1] ;
 wire \rvsingle.dp.rf.rf[13][20] ;
 wire \rvsingle.dp.rf.rf[13][21] ;
 wire \rvsingle.dp.rf.rf[13][22] ;
 wire \rvsingle.dp.rf.rf[13][23] ;
 wire \rvsingle.dp.rf.rf[13][24] ;
 wire \rvsingle.dp.rf.rf[13][25] ;
 wire \rvsingle.dp.rf.rf[13][26] ;
 wire \rvsingle.dp.rf.rf[13][27] ;
 wire \rvsingle.dp.rf.rf[13][28] ;
 wire \rvsingle.dp.rf.rf[13][29] ;
 wire \rvsingle.dp.rf.rf[13][2] ;
 wire \rvsingle.dp.rf.rf[13][30] ;
 wire \rvsingle.dp.rf.rf[13][31] ;
 wire \rvsingle.dp.rf.rf[13][3] ;
 wire \rvsingle.dp.rf.rf[13][4] ;
 wire \rvsingle.dp.rf.rf[13][5] ;
 wire \rvsingle.dp.rf.rf[13][6] ;
 wire \rvsingle.dp.rf.rf[13][7] ;
 wire \rvsingle.dp.rf.rf[13][8] ;
 wire \rvsingle.dp.rf.rf[13][9] ;
 wire \rvsingle.dp.rf.rf[14][0] ;
 wire \rvsingle.dp.rf.rf[14][10] ;
 wire \rvsingle.dp.rf.rf[14][11] ;
 wire \rvsingle.dp.rf.rf[14][12] ;
 wire \rvsingle.dp.rf.rf[14][13] ;
 wire \rvsingle.dp.rf.rf[14][14] ;
 wire \rvsingle.dp.rf.rf[14][15] ;
 wire \rvsingle.dp.rf.rf[14][16] ;
 wire \rvsingle.dp.rf.rf[14][17] ;
 wire \rvsingle.dp.rf.rf[14][18] ;
 wire \rvsingle.dp.rf.rf[14][19] ;
 wire \rvsingle.dp.rf.rf[14][1] ;
 wire \rvsingle.dp.rf.rf[14][20] ;
 wire \rvsingle.dp.rf.rf[14][21] ;
 wire \rvsingle.dp.rf.rf[14][22] ;
 wire \rvsingle.dp.rf.rf[14][23] ;
 wire \rvsingle.dp.rf.rf[14][24] ;
 wire \rvsingle.dp.rf.rf[14][25] ;
 wire \rvsingle.dp.rf.rf[14][26] ;
 wire \rvsingle.dp.rf.rf[14][27] ;
 wire \rvsingle.dp.rf.rf[14][28] ;
 wire \rvsingle.dp.rf.rf[14][29] ;
 wire \rvsingle.dp.rf.rf[14][2] ;
 wire \rvsingle.dp.rf.rf[14][30] ;
 wire \rvsingle.dp.rf.rf[14][31] ;
 wire \rvsingle.dp.rf.rf[14][3] ;
 wire \rvsingle.dp.rf.rf[14][4] ;
 wire \rvsingle.dp.rf.rf[14][5] ;
 wire \rvsingle.dp.rf.rf[14][6] ;
 wire \rvsingle.dp.rf.rf[14][7] ;
 wire \rvsingle.dp.rf.rf[14][8] ;
 wire \rvsingle.dp.rf.rf[14][9] ;
 wire \rvsingle.dp.rf.rf[15][0] ;
 wire \rvsingle.dp.rf.rf[15][10] ;
 wire \rvsingle.dp.rf.rf[15][11] ;
 wire \rvsingle.dp.rf.rf[15][12] ;
 wire \rvsingle.dp.rf.rf[15][13] ;
 wire \rvsingle.dp.rf.rf[15][14] ;
 wire \rvsingle.dp.rf.rf[15][15] ;
 wire \rvsingle.dp.rf.rf[15][16] ;
 wire \rvsingle.dp.rf.rf[15][17] ;
 wire \rvsingle.dp.rf.rf[15][18] ;
 wire \rvsingle.dp.rf.rf[15][19] ;
 wire \rvsingle.dp.rf.rf[15][1] ;
 wire \rvsingle.dp.rf.rf[15][20] ;
 wire \rvsingle.dp.rf.rf[15][21] ;
 wire \rvsingle.dp.rf.rf[15][22] ;
 wire \rvsingle.dp.rf.rf[15][23] ;
 wire \rvsingle.dp.rf.rf[15][24] ;
 wire \rvsingle.dp.rf.rf[15][25] ;
 wire \rvsingle.dp.rf.rf[15][26] ;
 wire \rvsingle.dp.rf.rf[15][27] ;
 wire \rvsingle.dp.rf.rf[15][28] ;
 wire \rvsingle.dp.rf.rf[15][29] ;
 wire \rvsingle.dp.rf.rf[15][2] ;
 wire \rvsingle.dp.rf.rf[15][30] ;
 wire \rvsingle.dp.rf.rf[15][31] ;
 wire \rvsingle.dp.rf.rf[15][3] ;
 wire \rvsingle.dp.rf.rf[15][4] ;
 wire \rvsingle.dp.rf.rf[15][5] ;
 wire \rvsingle.dp.rf.rf[15][6] ;
 wire \rvsingle.dp.rf.rf[15][7] ;
 wire \rvsingle.dp.rf.rf[15][8] ;
 wire \rvsingle.dp.rf.rf[15][9] ;
 wire \rvsingle.dp.rf.rf[16][0] ;
 wire \rvsingle.dp.rf.rf[16][10] ;
 wire \rvsingle.dp.rf.rf[16][11] ;
 wire \rvsingle.dp.rf.rf[16][12] ;
 wire \rvsingle.dp.rf.rf[16][13] ;
 wire \rvsingle.dp.rf.rf[16][14] ;
 wire \rvsingle.dp.rf.rf[16][15] ;
 wire \rvsingle.dp.rf.rf[16][16] ;
 wire \rvsingle.dp.rf.rf[16][17] ;
 wire \rvsingle.dp.rf.rf[16][18] ;
 wire \rvsingle.dp.rf.rf[16][19] ;
 wire \rvsingle.dp.rf.rf[16][1] ;
 wire \rvsingle.dp.rf.rf[16][20] ;
 wire \rvsingle.dp.rf.rf[16][21] ;
 wire \rvsingle.dp.rf.rf[16][22] ;
 wire \rvsingle.dp.rf.rf[16][23] ;
 wire \rvsingle.dp.rf.rf[16][24] ;
 wire \rvsingle.dp.rf.rf[16][25] ;
 wire \rvsingle.dp.rf.rf[16][26] ;
 wire \rvsingle.dp.rf.rf[16][27] ;
 wire \rvsingle.dp.rf.rf[16][28] ;
 wire \rvsingle.dp.rf.rf[16][29] ;
 wire \rvsingle.dp.rf.rf[16][2] ;
 wire \rvsingle.dp.rf.rf[16][30] ;
 wire \rvsingle.dp.rf.rf[16][31] ;
 wire \rvsingle.dp.rf.rf[16][3] ;
 wire \rvsingle.dp.rf.rf[16][4] ;
 wire \rvsingle.dp.rf.rf[16][5] ;
 wire \rvsingle.dp.rf.rf[16][6] ;
 wire \rvsingle.dp.rf.rf[16][7] ;
 wire \rvsingle.dp.rf.rf[16][8] ;
 wire \rvsingle.dp.rf.rf[16][9] ;
 wire \rvsingle.dp.rf.rf[17][0] ;
 wire \rvsingle.dp.rf.rf[17][10] ;
 wire \rvsingle.dp.rf.rf[17][11] ;
 wire \rvsingle.dp.rf.rf[17][12] ;
 wire \rvsingle.dp.rf.rf[17][13] ;
 wire \rvsingle.dp.rf.rf[17][14] ;
 wire \rvsingle.dp.rf.rf[17][15] ;
 wire \rvsingle.dp.rf.rf[17][16] ;
 wire \rvsingle.dp.rf.rf[17][17] ;
 wire \rvsingle.dp.rf.rf[17][18] ;
 wire \rvsingle.dp.rf.rf[17][19] ;
 wire \rvsingle.dp.rf.rf[17][1] ;
 wire \rvsingle.dp.rf.rf[17][20] ;
 wire \rvsingle.dp.rf.rf[17][21] ;
 wire \rvsingle.dp.rf.rf[17][22] ;
 wire \rvsingle.dp.rf.rf[17][23] ;
 wire \rvsingle.dp.rf.rf[17][24] ;
 wire \rvsingle.dp.rf.rf[17][25] ;
 wire \rvsingle.dp.rf.rf[17][26] ;
 wire \rvsingle.dp.rf.rf[17][27] ;
 wire \rvsingle.dp.rf.rf[17][28] ;
 wire \rvsingle.dp.rf.rf[17][29] ;
 wire \rvsingle.dp.rf.rf[17][2] ;
 wire \rvsingle.dp.rf.rf[17][30] ;
 wire \rvsingle.dp.rf.rf[17][31] ;
 wire \rvsingle.dp.rf.rf[17][3] ;
 wire \rvsingle.dp.rf.rf[17][4] ;
 wire \rvsingle.dp.rf.rf[17][5] ;
 wire \rvsingle.dp.rf.rf[17][6] ;
 wire \rvsingle.dp.rf.rf[17][7] ;
 wire \rvsingle.dp.rf.rf[17][8] ;
 wire \rvsingle.dp.rf.rf[17][9] ;
 wire \rvsingle.dp.rf.rf[18][0] ;
 wire \rvsingle.dp.rf.rf[18][10] ;
 wire \rvsingle.dp.rf.rf[18][11] ;
 wire \rvsingle.dp.rf.rf[18][12] ;
 wire \rvsingle.dp.rf.rf[18][13] ;
 wire \rvsingle.dp.rf.rf[18][14] ;
 wire \rvsingle.dp.rf.rf[18][15] ;
 wire \rvsingle.dp.rf.rf[18][16] ;
 wire \rvsingle.dp.rf.rf[18][17] ;
 wire \rvsingle.dp.rf.rf[18][18] ;
 wire \rvsingle.dp.rf.rf[18][19] ;
 wire \rvsingle.dp.rf.rf[18][1] ;
 wire \rvsingle.dp.rf.rf[18][20] ;
 wire \rvsingle.dp.rf.rf[18][21] ;
 wire \rvsingle.dp.rf.rf[18][22] ;
 wire \rvsingle.dp.rf.rf[18][23] ;
 wire \rvsingle.dp.rf.rf[18][24] ;
 wire \rvsingle.dp.rf.rf[18][25] ;
 wire \rvsingle.dp.rf.rf[18][26] ;
 wire \rvsingle.dp.rf.rf[18][27] ;
 wire \rvsingle.dp.rf.rf[18][28] ;
 wire \rvsingle.dp.rf.rf[18][29] ;
 wire \rvsingle.dp.rf.rf[18][2] ;
 wire \rvsingle.dp.rf.rf[18][30] ;
 wire \rvsingle.dp.rf.rf[18][31] ;
 wire \rvsingle.dp.rf.rf[18][3] ;
 wire \rvsingle.dp.rf.rf[18][4] ;
 wire \rvsingle.dp.rf.rf[18][5] ;
 wire \rvsingle.dp.rf.rf[18][6] ;
 wire \rvsingle.dp.rf.rf[18][7] ;
 wire \rvsingle.dp.rf.rf[18][8] ;
 wire \rvsingle.dp.rf.rf[18][9] ;
 wire \rvsingle.dp.rf.rf[19][0] ;
 wire \rvsingle.dp.rf.rf[19][10] ;
 wire \rvsingle.dp.rf.rf[19][11] ;
 wire \rvsingle.dp.rf.rf[19][12] ;
 wire \rvsingle.dp.rf.rf[19][13] ;
 wire \rvsingle.dp.rf.rf[19][14] ;
 wire \rvsingle.dp.rf.rf[19][15] ;
 wire \rvsingle.dp.rf.rf[19][16] ;
 wire \rvsingle.dp.rf.rf[19][17] ;
 wire \rvsingle.dp.rf.rf[19][18] ;
 wire \rvsingle.dp.rf.rf[19][19] ;
 wire \rvsingle.dp.rf.rf[19][1] ;
 wire \rvsingle.dp.rf.rf[19][20] ;
 wire \rvsingle.dp.rf.rf[19][21] ;
 wire \rvsingle.dp.rf.rf[19][22] ;
 wire \rvsingle.dp.rf.rf[19][23] ;
 wire \rvsingle.dp.rf.rf[19][24] ;
 wire \rvsingle.dp.rf.rf[19][25] ;
 wire \rvsingle.dp.rf.rf[19][26] ;
 wire \rvsingle.dp.rf.rf[19][27] ;
 wire \rvsingle.dp.rf.rf[19][28] ;
 wire \rvsingle.dp.rf.rf[19][29] ;
 wire \rvsingle.dp.rf.rf[19][2] ;
 wire \rvsingle.dp.rf.rf[19][30] ;
 wire \rvsingle.dp.rf.rf[19][31] ;
 wire \rvsingle.dp.rf.rf[19][3] ;
 wire \rvsingle.dp.rf.rf[19][4] ;
 wire \rvsingle.dp.rf.rf[19][5] ;
 wire \rvsingle.dp.rf.rf[19][6] ;
 wire \rvsingle.dp.rf.rf[19][7] ;
 wire \rvsingle.dp.rf.rf[19][8] ;
 wire \rvsingle.dp.rf.rf[19][9] ;
 wire \rvsingle.dp.rf.rf[1][0] ;
 wire \rvsingle.dp.rf.rf[1][10] ;
 wire \rvsingle.dp.rf.rf[1][11] ;
 wire \rvsingle.dp.rf.rf[1][12] ;
 wire \rvsingle.dp.rf.rf[1][13] ;
 wire \rvsingle.dp.rf.rf[1][14] ;
 wire \rvsingle.dp.rf.rf[1][15] ;
 wire \rvsingle.dp.rf.rf[1][16] ;
 wire \rvsingle.dp.rf.rf[1][17] ;
 wire \rvsingle.dp.rf.rf[1][18] ;
 wire \rvsingle.dp.rf.rf[1][19] ;
 wire \rvsingle.dp.rf.rf[1][1] ;
 wire \rvsingle.dp.rf.rf[1][20] ;
 wire \rvsingle.dp.rf.rf[1][21] ;
 wire \rvsingle.dp.rf.rf[1][22] ;
 wire \rvsingle.dp.rf.rf[1][23] ;
 wire \rvsingle.dp.rf.rf[1][24] ;
 wire \rvsingle.dp.rf.rf[1][25] ;
 wire \rvsingle.dp.rf.rf[1][26] ;
 wire \rvsingle.dp.rf.rf[1][27] ;
 wire \rvsingle.dp.rf.rf[1][28] ;
 wire \rvsingle.dp.rf.rf[1][29] ;
 wire \rvsingle.dp.rf.rf[1][2] ;
 wire \rvsingle.dp.rf.rf[1][30] ;
 wire \rvsingle.dp.rf.rf[1][31] ;
 wire \rvsingle.dp.rf.rf[1][3] ;
 wire \rvsingle.dp.rf.rf[1][4] ;
 wire \rvsingle.dp.rf.rf[1][5] ;
 wire \rvsingle.dp.rf.rf[1][6] ;
 wire \rvsingle.dp.rf.rf[1][7] ;
 wire \rvsingle.dp.rf.rf[1][8] ;
 wire \rvsingle.dp.rf.rf[1][9] ;
 wire \rvsingle.dp.rf.rf[20][0] ;
 wire \rvsingle.dp.rf.rf[20][10] ;
 wire \rvsingle.dp.rf.rf[20][11] ;
 wire \rvsingle.dp.rf.rf[20][12] ;
 wire \rvsingle.dp.rf.rf[20][13] ;
 wire \rvsingle.dp.rf.rf[20][14] ;
 wire \rvsingle.dp.rf.rf[20][15] ;
 wire \rvsingle.dp.rf.rf[20][16] ;
 wire \rvsingle.dp.rf.rf[20][17] ;
 wire \rvsingle.dp.rf.rf[20][18] ;
 wire \rvsingle.dp.rf.rf[20][19] ;
 wire \rvsingle.dp.rf.rf[20][1] ;
 wire \rvsingle.dp.rf.rf[20][20] ;
 wire \rvsingle.dp.rf.rf[20][21] ;
 wire \rvsingle.dp.rf.rf[20][22] ;
 wire \rvsingle.dp.rf.rf[20][23] ;
 wire \rvsingle.dp.rf.rf[20][24] ;
 wire \rvsingle.dp.rf.rf[20][25] ;
 wire \rvsingle.dp.rf.rf[20][26] ;
 wire \rvsingle.dp.rf.rf[20][27] ;
 wire \rvsingle.dp.rf.rf[20][28] ;
 wire \rvsingle.dp.rf.rf[20][29] ;
 wire \rvsingle.dp.rf.rf[20][2] ;
 wire \rvsingle.dp.rf.rf[20][30] ;
 wire \rvsingle.dp.rf.rf[20][31] ;
 wire \rvsingle.dp.rf.rf[20][3] ;
 wire \rvsingle.dp.rf.rf[20][4] ;
 wire \rvsingle.dp.rf.rf[20][5] ;
 wire \rvsingle.dp.rf.rf[20][6] ;
 wire \rvsingle.dp.rf.rf[20][7] ;
 wire \rvsingle.dp.rf.rf[20][8] ;
 wire \rvsingle.dp.rf.rf[20][9] ;
 wire \rvsingle.dp.rf.rf[21][0] ;
 wire \rvsingle.dp.rf.rf[21][10] ;
 wire \rvsingle.dp.rf.rf[21][11] ;
 wire \rvsingle.dp.rf.rf[21][12] ;
 wire \rvsingle.dp.rf.rf[21][13] ;
 wire \rvsingle.dp.rf.rf[21][14] ;
 wire \rvsingle.dp.rf.rf[21][15] ;
 wire \rvsingle.dp.rf.rf[21][16] ;
 wire \rvsingle.dp.rf.rf[21][17] ;
 wire \rvsingle.dp.rf.rf[21][18] ;
 wire \rvsingle.dp.rf.rf[21][19] ;
 wire \rvsingle.dp.rf.rf[21][1] ;
 wire \rvsingle.dp.rf.rf[21][20] ;
 wire \rvsingle.dp.rf.rf[21][21] ;
 wire \rvsingle.dp.rf.rf[21][22] ;
 wire \rvsingle.dp.rf.rf[21][23] ;
 wire \rvsingle.dp.rf.rf[21][24] ;
 wire \rvsingle.dp.rf.rf[21][25] ;
 wire \rvsingle.dp.rf.rf[21][26] ;
 wire \rvsingle.dp.rf.rf[21][27] ;
 wire \rvsingle.dp.rf.rf[21][28] ;
 wire \rvsingle.dp.rf.rf[21][29] ;
 wire \rvsingle.dp.rf.rf[21][2] ;
 wire \rvsingle.dp.rf.rf[21][30] ;
 wire \rvsingle.dp.rf.rf[21][31] ;
 wire \rvsingle.dp.rf.rf[21][3] ;
 wire \rvsingle.dp.rf.rf[21][4] ;
 wire \rvsingle.dp.rf.rf[21][5] ;
 wire \rvsingle.dp.rf.rf[21][6] ;
 wire \rvsingle.dp.rf.rf[21][7] ;
 wire \rvsingle.dp.rf.rf[21][8] ;
 wire \rvsingle.dp.rf.rf[21][9] ;
 wire \rvsingle.dp.rf.rf[22][0] ;
 wire \rvsingle.dp.rf.rf[22][10] ;
 wire \rvsingle.dp.rf.rf[22][11] ;
 wire \rvsingle.dp.rf.rf[22][12] ;
 wire \rvsingle.dp.rf.rf[22][13] ;
 wire \rvsingle.dp.rf.rf[22][14] ;
 wire \rvsingle.dp.rf.rf[22][15] ;
 wire \rvsingle.dp.rf.rf[22][16] ;
 wire \rvsingle.dp.rf.rf[22][17] ;
 wire \rvsingle.dp.rf.rf[22][18] ;
 wire \rvsingle.dp.rf.rf[22][19] ;
 wire \rvsingle.dp.rf.rf[22][1] ;
 wire \rvsingle.dp.rf.rf[22][20] ;
 wire \rvsingle.dp.rf.rf[22][21] ;
 wire \rvsingle.dp.rf.rf[22][22] ;
 wire \rvsingle.dp.rf.rf[22][23] ;
 wire \rvsingle.dp.rf.rf[22][24] ;
 wire \rvsingle.dp.rf.rf[22][25] ;
 wire \rvsingle.dp.rf.rf[22][26] ;
 wire \rvsingle.dp.rf.rf[22][27] ;
 wire \rvsingle.dp.rf.rf[22][28] ;
 wire \rvsingle.dp.rf.rf[22][29] ;
 wire \rvsingle.dp.rf.rf[22][2] ;
 wire \rvsingle.dp.rf.rf[22][30] ;
 wire \rvsingle.dp.rf.rf[22][31] ;
 wire \rvsingle.dp.rf.rf[22][3] ;
 wire \rvsingle.dp.rf.rf[22][4] ;
 wire \rvsingle.dp.rf.rf[22][5] ;
 wire \rvsingle.dp.rf.rf[22][6] ;
 wire \rvsingle.dp.rf.rf[22][7] ;
 wire \rvsingle.dp.rf.rf[22][8] ;
 wire \rvsingle.dp.rf.rf[22][9] ;
 wire \rvsingle.dp.rf.rf[23][0] ;
 wire \rvsingle.dp.rf.rf[23][10] ;
 wire \rvsingle.dp.rf.rf[23][11] ;
 wire \rvsingle.dp.rf.rf[23][12] ;
 wire \rvsingle.dp.rf.rf[23][13] ;
 wire \rvsingle.dp.rf.rf[23][14] ;
 wire \rvsingle.dp.rf.rf[23][15] ;
 wire \rvsingle.dp.rf.rf[23][16] ;
 wire \rvsingle.dp.rf.rf[23][17] ;
 wire \rvsingle.dp.rf.rf[23][18] ;
 wire \rvsingle.dp.rf.rf[23][19] ;
 wire \rvsingle.dp.rf.rf[23][1] ;
 wire \rvsingle.dp.rf.rf[23][20] ;
 wire \rvsingle.dp.rf.rf[23][21] ;
 wire \rvsingle.dp.rf.rf[23][22] ;
 wire \rvsingle.dp.rf.rf[23][23] ;
 wire \rvsingle.dp.rf.rf[23][24] ;
 wire \rvsingle.dp.rf.rf[23][25] ;
 wire \rvsingle.dp.rf.rf[23][26] ;
 wire \rvsingle.dp.rf.rf[23][27] ;
 wire \rvsingle.dp.rf.rf[23][28] ;
 wire \rvsingle.dp.rf.rf[23][29] ;
 wire \rvsingle.dp.rf.rf[23][2] ;
 wire \rvsingle.dp.rf.rf[23][30] ;
 wire \rvsingle.dp.rf.rf[23][31] ;
 wire \rvsingle.dp.rf.rf[23][3] ;
 wire \rvsingle.dp.rf.rf[23][4] ;
 wire \rvsingle.dp.rf.rf[23][5] ;
 wire \rvsingle.dp.rf.rf[23][6] ;
 wire \rvsingle.dp.rf.rf[23][7] ;
 wire \rvsingle.dp.rf.rf[23][8] ;
 wire \rvsingle.dp.rf.rf[23][9] ;
 wire \rvsingle.dp.rf.rf[24][0] ;
 wire \rvsingle.dp.rf.rf[24][10] ;
 wire \rvsingle.dp.rf.rf[24][11] ;
 wire \rvsingle.dp.rf.rf[24][12] ;
 wire \rvsingle.dp.rf.rf[24][13] ;
 wire \rvsingle.dp.rf.rf[24][14] ;
 wire \rvsingle.dp.rf.rf[24][15] ;
 wire \rvsingle.dp.rf.rf[24][16] ;
 wire \rvsingle.dp.rf.rf[24][17] ;
 wire \rvsingle.dp.rf.rf[24][18] ;
 wire \rvsingle.dp.rf.rf[24][19] ;
 wire \rvsingle.dp.rf.rf[24][1] ;
 wire \rvsingle.dp.rf.rf[24][20] ;
 wire \rvsingle.dp.rf.rf[24][21] ;
 wire \rvsingle.dp.rf.rf[24][22] ;
 wire \rvsingle.dp.rf.rf[24][23] ;
 wire \rvsingle.dp.rf.rf[24][24] ;
 wire \rvsingle.dp.rf.rf[24][25] ;
 wire \rvsingle.dp.rf.rf[24][26] ;
 wire \rvsingle.dp.rf.rf[24][27] ;
 wire \rvsingle.dp.rf.rf[24][28] ;
 wire \rvsingle.dp.rf.rf[24][29] ;
 wire \rvsingle.dp.rf.rf[24][2] ;
 wire \rvsingle.dp.rf.rf[24][30] ;
 wire \rvsingle.dp.rf.rf[24][31] ;
 wire \rvsingle.dp.rf.rf[24][3] ;
 wire \rvsingle.dp.rf.rf[24][4] ;
 wire \rvsingle.dp.rf.rf[24][5] ;
 wire \rvsingle.dp.rf.rf[24][6] ;
 wire \rvsingle.dp.rf.rf[24][7] ;
 wire \rvsingle.dp.rf.rf[24][8] ;
 wire \rvsingle.dp.rf.rf[24][9] ;
 wire \rvsingle.dp.rf.rf[25][0] ;
 wire \rvsingle.dp.rf.rf[25][10] ;
 wire \rvsingle.dp.rf.rf[25][11] ;
 wire \rvsingle.dp.rf.rf[25][12] ;
 wire \rvsingle.dp.rf.rf[25][13] ;
 wire \rvsingle.dp.rf.rf[25][14] ;
 wire \rvsingle.dp.rf.rf[25][15] ;
 wire \rvsingle.dp.rf.rf[25][16] ;
 wire \rvsingle.dp.rf.rf[25][17] ;
 wire \rvsingle.dp.rf.rf[25][18] ;
 wire \rvsingle.dp.rf.rf[25][19] ;
 wire \rvsingle.dp.rf.rf[25][1] ;
 wire \rvsingle.dp.rf.rf[25][20] ;
 wire \rvsingle.dp.rf.rf[25][21] ;
 wire \rvsingle.dp.rf.rf[25][22] ;
 wire \rvsingle.dp.rf.rf[25][23] ;
 wire \rvsingle.dp.rf.rf[25][24] ;
 wire \rvsingle.dp.rf.rf[25][25] ;
 wire \rvsingle.dp.rf.rf[25][26] ;
 wire \rvsingle.dp.rf.rf[25][27] ;
 wire \rvsingle.dp.rf.rf[25][28] ;
 wire \rvsingle.dp.rf.rf[25][29] ;
 wire \rvsingle.dp.rf.rf[25][2] ;
 wire \rvsingle.dp.rf.rf[25][30] ;
 wire \rvsingle.dp.rf.rf[25][31] ;
 wire \rvsingle.dp.rf.rf[25][3] ;
 wire \rvsingle.dp.rf.rf[25][4] ;
 wire \rvsingle.dp.rf.rf[25][5] ;
 wire \rvsingle.dp.rf.rf[25][6] ;
 wire \rvsingle.dp.rf.rf[25][7] ;
 wire \rvsingle.dp.rf.rf[25][8] ;
 wire \rvsingle.dp.rf.rf[25][9] ;
 wire \rvsingle.dp.rf.rf[26][0] ;
 wire \rvsingle.dp.rf.rf[26][10] ;
 wire \rvsingle.dp.rf.rf[26][11] ;
 wire \rvsingle.dp.rf.rf[26][12] ;
 wire \rvsingle.dp.rf.rf[26][13] ;
 wire \rvsingle.dp.rf.rf[26][14] ;
 wire \rvsingle.dp.rf.rf[26][15] ;
 wire \rvsingle.dp.rf.rf[26][16] ;
 wire \rvsingle.dp.rf.rf[26][17] ;
 wire \rvsingle.dp.rf.rf[26][18] ;
 wire \rvsingle.dp.rf.rf[26][19] ;
 wire \rvsingle.dp.rf.rf[26][1] ;
 wire \rvsingle.dp.rf.rf[26][20] ;
 wire \rvsingle.dp.rf.rf[26][21] ;
 wire \rvsingle.dp.rf.rf[26][22] ;
 wire \rvsingle.dp.rf.rf[26][23] ;
 wire \rvsingle.dp.rf.rf[26][24] ;
 wire \rvsingle.dp.rf.rf[26][25] ;
 wire \rvsingle.dp.rf.rf[26][26] ;
 wire \rvsingle.dp.rf.rf[26][27] ;
 wire \rvsingle.dp.rf.rf[26][28] ;
 wire \rvsingle.dp.rf.rf[26][29] ;
 wire \rvsingle.dp.rf.rf[26][2] ;
 wire \rvsingle.dp.rf.rf[26][30] ;
 wire \rvsingle.dp.rf.rf[26][31] ;
 wire \rvsingle.dp.rf.rf[26][3] ;
 wire \rvsingle.dp.rf.rf[26][4] ;
 wire \rvsingle.dp.rf.rf[26][5] ;
 wire \rvsingle.dp.rf.rf[26][6] ;
 wire \rvsingle.dp.rf.rf[26][7] ;
 wire \rvsingle.dp.rf.rf[26][8] ;
 wire \rvsingle.dp.rf.rf[26][9] ;
 wire \rvsingle.dp.rf.rf[27][0] ;
 wire \rvsingle.dp.rf.rf[27][10] ;
 wire \rvsingle.dp.rf.rf[27][11] ;
 wire \rvsingle.dp.rf.rf[27][12] ;
 wire \rvsingle.dp.rf.rf[27][13] ;
 wire \rvsingle.dp.rf.rf[27][14] ;
 wire \rvsingle.dp.rf.rf[27][15] ;
 wire \rvsingle.dp.rf.rf[27][16] ;
 wire \rvsingle.dp.rf.rf[27][17] ;
 wire \rvsingle.dp.rf.rf[27][18] ;
 wire \rvsingle.dp.rf.rf[27][19] ;
 wire \rvsingle.dp.rf.rf[27][1] ;
 wire \rvsingle.dp.rf.rf[27][20] ;
 wire \rvsingle.dp.rf.rf[27][21] ;
 wire \rvsingle.dp.rf.rf[27][22] ;
 wire \rvsingle.dp.rf.rf[27][23] ;
 wire \rvsingle.dp.rf.rf[27][24] ;
 wire \rvsingle.dp.rf.rf[27][25] ;
 wire \rvsingle.dp.rf.rf[27][26] ;
 wire \rvsingle.dp.rf.rf[27][27] ;
 wire \rvsingle.dp.rf.rf[27][28] ;
 wire \rvsingle.dp.rf.rf[27][29] ;
 wire \rvsingle.dp.rf.rf[27][2] ;
 wire \rvsingle.dp.rf.rf[27][30] ;
 wire \rvsingle.dp.rf.rf[27][31] ;
 wire \rvsingle.dp.rf.rf[27][3] ;
 wire \rvsingle.dp.rf.rf[27][4] ;
 wire \rvsingle.dp.rf.rf[27][5] ;
 wire \rvsingle.dp.rf.rf[27][6] ;
 wire \rvsingle.dp.rf.rf[27][7] ;
 wire \rvsingle.dp.rf.rf[27][8] ;
 wire \rvsingle.dp.rf.rf[27][9] ;
 wire \rvsingle.dp.rf.rf[28][0] ;
 wire \rvsingle.dp.rf.rf[28][10] ;
 wire \rvsingle.dp.rf.rf[28][11] ;
 wire \rvsingle.dp.rf.rf[28][12] ;
 wire \rvsingle.dp.rf.rf[28][13] ;
 wire \rvsingle.dp.rf.rf[28][14] ;
 wire \rvsingle.dp.rf.rf[28][15] ;
 wire \rvsingle.dp.rf.rf[28][16] ;
 wire \rvsingle.dp.rf.rf[28][17] ;
 wire \rvsingle.dp.rf.rf[28][18] ;
 wire \rvsingle.dp.rf.rf[28][19] ;
 wire \rvsingle.dp.rf.rf[28][1] ;
 wire \rvsingle.dp.rf.rf[28][20] ;
 wire \rvsingle.dp.rf.rf[28][21] ;
 wire \rvsingle.dp.rf.rf[28][22] ;
 wire \rvsingle.dp.rf.rf[28][23] ;
 wire \rvsingle.dp.rf.rf[28][24] ;
 wire \rvsingle.dp.rf.rf[28][25] ;
 wire \rvsingle.dp.rf.rf[28][26] ;
 wire \rvsingle.dp.rf.rf[28][27] ;
 wire \rvsingle.dp.rf.rf[28][28] ;
 wire \rvsingle.dp.rf.rf[28][29] ;
 wire \rvsingle.dp.rf.rf[28][2] ;
 wire \rvsingle.dp.rf.rf[28][30] ;
 wire \rvsingle.dp.rf.rf[28][31] ;
 wire \rvsingle.dp.rf.rf[28][3] ;
 wire \rvsingle.dp.rf.rf[28][4] ;
 wire \rvsingle.dp.rf.rf[28][5] ;
 wire \rvsingle.dp.rf.rf[28][6] ;
 wire \rvsingle.dp.rf.rf[28][7] ;
 wire \rvsingle.dp.rf.rf[28][8] ;
 wire \rvsingle.dp.rf.rf[28][9] ;
 wire \rvsingle.dp.rf.rf[29][0] ;
 wire \rvsingle.dp.rf.rf[29][10] ;
 wire \rvsingle.dp.rf.rf[29][11] ;
 wire \rvsingle.dp.rf.rf[29][12] ;
 wire \rvsingle.dp.rf.rf[29][13] ;
 wire \rvsingle.dp.rf.rf[29][14] ;
 wire \rvsingle.dp.rf.rf[29][15] ;
 wire \rvsingle.dp.rf.rf[29][16] ;
 wire \rvsingle.dp.rf.rf[29][17] ;
 wire \rvsingle.dp.rf.rf[29][18] ;
 wire \rvsingle.dp.rf.rf[29][19] ;
 wire \rvsingle.dp.rf.rf[29][1] ;
 wire \rvsingle.dp.rf.rf[29][20] ;
 wire \rvsingle.dp.rf.rf[29][21] ;
 wire \rvsingle.dp.rf.rf[29][22] ;
 wire \rvsingle.dp.rf.rf[29][23] ;
 wire \rvsingle.dp.rf.rf[29][24] ;
 wire \rvsingle.dp.rf.rf[29][25] ;
 wire \rvsingle.dp.rf.rf[29][26] ;
 wire \rvsingle.dp.rf.rf[29][27] ;
 wire \rvsingle.dp.rf.rf[29][28] ;
 wire \rvsingle.dp.rf.rf[29][29] ;
 wire \rvsingle.dp.rf.rf[29][2] ;
 wire \rvsingle.dp.rf.rf[29][30] ;
 wire \rvsingle.dp.rf.rf[29][31] ;
 wire \rvsingle.dp.rf.rf[29][3] ;
 wire \rvsingle.dp.rf.rf[29][4] ;
 wire \rvsingle.dp.rf.rf[29][5] ;
 wire \rvsingle.dp.rf.rf[29][6] ;
 wire \rvsingle.dp.rf.rf[29][7] ;
 wire \rvsingle.dp.rf.rf[29][8] ;
 wire \rvsingle.dp.rf.rf[29][9] ;
 wire \rvsingle.dp.rf.rf[2][0] ;
 wire \rvsingle.dp.rf.rf[2][10] ;
 wire \rvsingle.dp.rf.rf[2][11] ;
 wire \rvsingle.dp.rf.rf[2][12] ;
 wire \rvsingle.dp.rf.rf[2][13] ;
 wire \rvsingle.dp.rf.rf[2][14] ;
 wire \rvsingle.dp.rf.rf[2][15] ;
 wire \rvsingle.dp.rf.rf[2][16] ;
 wire \rvsingle.dp.rf.rf[2][17] ;
 wire \rvsingle.dp.rf.rf[2][18] ;
 wire \rvsingle.dp.rf.rf[2][19] ;
 wire \rvsingle.dp.rf.rf[2][1] ;
 wire \rvsingle.dp.rf.rf[2][20] ;
 wire \rvsingle.dp.rf.rf[2][21] ;
 wire \rvsingle.dp.rf.rf[2][22] ;
 wire \rvsingle.dp.rf.rf[2][23] ;
 wire \rvsingle.dp.rf.rf[2][24] ;
 wire \rvsingle.dp.rf.rf[2][25] ;
 wire \rvsingle.dp.rf.rf[2][26] ;
 wire \rvsingle.dp.rf.rf[2][27] ;
 wire \rvsingle.dp.rf.rf[2][28] ;
 wire \rvsingle.dp.rf.rf[2][29] ;
 wire \rvsingle.dp.rf.rf[2][2] ;
 wire \rvsingle.dp.rf.rf[2][30] ;
 wire \rvsingle.dp.rf.rf[2][31] ;
 wire \rvsingle.dp.rf.rf[2][3] ;
 wire \rvsingle.dp.rf.rf[2][4] ;
 wire \rvsingle.dp.rf.rf[2][5] ;
 wire \rvsingle.dp.rf.rf[2][6] ;
 wire \rvsingle.dp.rf.rf[2][7] ;
 wire \rvsingle.dp.rf.rf[2][8] ;
 wire \rvsingle.dp.rf.rf[2][9] ;
 wire \rvsingle.dp.rf.rf[30][0] ;
 wire \rvsingle.dp.rf.rf[30][10] ;
 wire \rvsingle.dp.rf.rf[30][11] ;
 wire \rvsingle.dp.rf.rf[30][12] ;
 wire \rvsingle.dp.rf.rf[30][13] ;
 wire \rvsingle.dp.rf.rf[30][14] ;
 wire \rvsingle.dp.rf.rf[30][15] ;
 wire \rvsingle.dp.rf.rf[30][16] ;
 wire \rvsingle.dp.rf.rf[30][17] ;
 wire \rvsingle.dp.rf.rf[30][18] ;
 wire \rvsingle.dp.rf.rf[30][19] ;
 wire \rvsingle.dp.rf.rf[30][1] ;
 wire \rvsingle.dp.rf.rf[30][20] ;
 wire \rvsingle.dp.rf.rf[30][21] ;
 wire \rvsingle.dp.rf.rf[30][22] ;
 wire \rvsingle.dp.rf.rf[30][23] ;
 wire \rvsingle.dp.rf.rf[30][24] ;
 wire \rvsingle.dp.rf.rf[30][25] ;
 wire \rvsingle.dp.rf.rf[30][26] ;
 wire \rvsingle.dp.rf.rf[30][27] ;
 wire \rvsingle.dp.rf.rf[30][28] ;
 wire \rvsingle.dp.rf.rf[30][29] ;
 wire \rvsingle.dp.rf.rf[30][2] ;
 wire \rvsingle.dp.rf.rf[30][30] ;
 wire \rvsingle.dp.rf.rf[30][31] ;
 wire \rvsingle.dp.rf.rf[30][3] ;
 wire \rvsingle.dp.rf.rf[30][4] ;
 wire \rvsingle.dp.rf.rf[30][5] ;
 wire \rvsingle.dp.rf.rf[30][6] ;
 wire \rvsingle.dp.rf.rf[30][7] ;
 wire \rvsingle.dp.rf.rf[30][8] ;
 wire \rvsingle.dp.rf.rf[30][9] ;
 wire \rvsingle.dp.rf.rf[31][0] ;
 wire \rvsingle.dp.rf.rf[31][10] ;
 wire \rvsingle.dp.rf.rf[31][11] ;
 wire \rvsingle.dp.rf.rf[31][12] ;
 wire \rvsingle.dp.rf.rf[31][13] ;
 wire \rvsingle.dp.rf.rf[31][14] ;
 wire \rvsingle.dp.rf.rf[31][15] ;
 wire \rvsingle.dp.rf.rf[31][16] ;
 wire \rvsingle.dp.rf.rf[31][17] ;
 wire \rvsingle.dp.rf.rf[31][18] ;
 wire \rvsingle.dp.rf.rf[31][19] ;
 wire \rvsingle.dp.rf.rf[31][1] ;
 wire \rvsingle.dp.rf.rf[31][20] ;
 wire \rvsingle.dp.rf.rf[31][21] ;
 wire \rvsingle.dp.rf.rf[31][22] ;
 wire \rvsingle.dp.rf.rf[31][23] ;
 wire \rvsingle.dp.rf.rf[31][24] ;
 wire \rvsingle.dp.rf.rf[31][25] ;
 wire \rvsingle.dp.rf.rf[31][26] ;
 wire \rvsingle.dp.rf.rf[31][27] ;
 wire \rvsingle.dp.rf.rf[31][28] ;
 wire \rvsingle.dp.rf.rf[31][29] ;
 wire \rvsingle.dp.rf.rf[31][2] ;
 wire \rvsingle.dp.rf.rf[31][30] ;
 wire \rvsingle.dp.rf.rf[31][31] ;
 wire \rvsingle.dp.rf.rf[31][3] ;
 wire \rvsingle.dp.rf.rf[31][4] ;
 wire \rvsingle.dp.rf.rf[31][5] ;
 wire \rvsingle.dp.rf.rf[31][6] ;
 wire \rvsingle.dp.rf.rf[31][7] ;
 wire \rvsingle.dp.rf.rf[31][8] ;
 wire \rvsingle.dp.rf.rf[31][9] ;
 wire \rvsingle.dp.rf.rf[3][0] ;
 wire \rvsingle.dp.rf.rf[3][10] ;
 wire \rvsingle.dp.rf.rf[3][11] ;
 wire \rvsingle.dp.rf.rf[3][12] ;
 wire \rvsingle.dp.rf.rf[3][13] ;
 wire \rvsingle.dp.rf.rf[3][14] ;
 wire \rvsingle.dp.rf.rf[3][15] ;
 wire \rvsingle.dp.rf.rf[3][16] ;
 wire \rvsingle.dp.rf.rf[3][17] ;
 wire \rvsingle.dp.rf.rf[3][18] ;
 wire \rvsingle.dp.rf.rf[3][19] ;
 wire \rvsingle.dp.rf.rf[3][1] ;
 wire \rvsingle.dp.rf.rf[3][20] ;
 wire \rvsingle.dp.rf.rf[3][21] ;
 wire \rvsingle.dp.rf.rf[3][22] ;
 wire \rvsingle.dp.rf.rf[3][23] ;
 wire \rvsingle.dp.rf.rf[3][24] ;
 wire \rvsingle.dp.rf.rf[3][25] ;
 wire \rvsingle.dp.rf.rf[3][26] ;
 wire \rvsingle.dp.rf.rf[3][27] ;
 wire \rvsingle.dp.rf.rf[3][28] ;
 wire \rvsingle.dp.rf.rf[3][29] ;
 wire \rvsingle.dp.rf.rf[3][2] ;
 wire \rvsingle.dp.rf.rf[3][30] ;
 wire \rvsingle.dp.rf.rf[3][31] ;
 wire \rvsingle.dp.rf.rf[3][3] ;
 wire \rvsingle.dp.rf.rf[3][4] ;
 wire \rvsingle.dp.rf.rf[3][5] ;
 wire \rvsingle.dp.rf.rf[3][6] ;
 wire \rvsingle.dp.rf.rf[3][7] ;
 wire \rvsingle.dp.rf.rf[3][8] ;
 wire \rvsingle.dp.rf.rf[3][9] ;
 wire \rvsingle.dp.rf.rf[4][0] ;
 wire \rvsingle.dp.rf.rf[4][10] ;
 wire \rvsingle.dp.rf.rf[4][11] ;
 wire \rvsingle.dp.rf.rf[4][12] ;
 wire \rvsingle.dp.rf.rf[4][13] ;
 wire \rvsingle.dp.rf.rf[4][14] ;
 wire \rvsingle.dp.rf.rf[4][15] ;
 wire \rvsingle.dp.rf.rf[4][16] ;
 wire \rvsingle.dp.rf.rf[4][17] ;
 wire \rvsingle.dp.rf.rf[4][18] ;
 wire \rvsingle.dp.rf.rf[4][19] ;
 wire \rvsingle.dp.rf.rf[4][1] ;
 wire \rvsingle.dp.rf.rf[4][20] ;
 wire \rvsingle.dp.rf.rf[4][21] ;
 wire \rvsingle.dp.rf.rf[4][22] ;
 wire \rvsingle.dp.rf.rf[4][23] ;
 wire \rvsingle.dp.rf.rf[4][24] ;
 wire \rvsingle.dp.rf.rf[4][25] ;
 wire \rvsingle.dp.rf.rf[4][26] ;
 wire \rvsingle.dp.rf.rf[4][27] ;
 wire \rvsingle.dp.rf.rf[4][28] ;
 wire \rvsingle.dp.rf.rf[4][29] ;
 wire \rvsingle.dp.rf.rf[4][2] ;
 wire \rvsingle.dp.rf.rf[4][30] ;
 wire \rvsingle.dp.rf.rf[4][31] ;
 wire \rvsingle.dp.rf.rf[4][3] ;
 wire \rvsingle.dp.rf.rf[4][4] ;
 wire \rvsingle.dp.rf.rf[4][5] ;
 wire \rvsingle.dp.rf.rf[4][6] ;
 wire \rvsingle.dp.rf.rf[4][7] ;
 wire \rvsingle.dp.rf.rf[4][8] ;
 wire \rvsingle.dp.rf.rf[4][9] ;
 wire \rvsingle.dp.rf.rf[5][0] ;
 wire \rvsingle.dp.rf.rf[5][10] ;
 wire \rvsingle.dp.rf.rf[5][11] ;
 wire \rvsingle.dp.rf.rf[5][12] ;
 wire \rvsingle.dp.rf.rf[5][13] ;
 wire \rvsingle.dp.rf.rf[5][14] ;
 wire \rvsingle.dp.rf.rf[5][15] ;
 wire \rvsingle.dp.rf.rf[5][16] ;
 wire \rvsingle.dp.rf.rf[5][17] ;
 wire \rvsingle.dp.rf.rf[5][18] ;
 wire \rvsingle.dp.rf.rf[5][19] ;
 wire \rvsingle.dp.rf.rf[5][1] ;
 wire \rvsingle.dp.rf.rf[5][20] ;
 wire \rvsingle.dp.rf.rf[5][21] ;
 wire \rvsingle.dp.rf.rf[5][22] ;
 wire \rvsingle.dp.rf.rf[5][23] ;
 wire \rvsingle.dp.rf.rf[5][24] ;
 wire \rvsingle.dp.rf.rf[5][25] ;
 wire \rvsingle.dp.rf.rf[5][26] ;
 wire \rvsingle.dp.rf.rf[5][27] ;
 wire \rvsingle.dp.rf.rf[5][28] ;
 wire \rvsingle.dp.rf.rf[5][29] ;
 wire \rvsingle.dp.rf.rf[5][2] ;
 wire \rvsingle.dp.rf.rf[5][30] ;
 wire \rvsingle.dp.rf.rf[5][31] ;
 wire \rvsingle.dp.rf.rf[5][3] ;
 wire \rvsingle.dp.rf.rf[5][4] ;
 wire \rvsingle.dp.rf.rf[5][5] ;
 wire \rvsingle.dp.rf.rf[5][6] ;
 wire \rvsingle.dp.rf.rf[5][7] ;
 wire \rvsingle.dp.rf.rf[5][8] ;
 wire \rvsingle.dp.rf.rf[5][9] ;
 wire \rvsingle.dp.rf.rf[6][0] ;
 wire \rvsingle.dp.rf.rf[6][10] ;
 wire \rvsingle.dp.rf.rf[6][11] ;
 wire \rvsingle.dp.rf.rf[6][12] ;
 wire \rvsingle.dp.rf.rf[6][13] ;
 wire \rvsingle.dp.rf.rf[6][14] ;
 wire \rvsingle.dp.rf.rf[6][15] ;
 wire \rvsingle.dp.rf.rf[6][16] ;
 wire \rvsingle.dp.rf.rf[6][17] ;
 wire \rvsingle.dp.rf.rf[6][18] ;
 wire \rvsingle.dp.rf.rf[6][19] ;
 wire \rvsingle.dp.rf.rf[6][1] ;
 wire \rvsingle.dp.rf.rf[6][20] ;
 wire \rvsingle.dp.rf.rf[6][21] ;
 wire \rvsingle.dp.rf.rf[6][22] ;
 wire \rvsingle.dp.rf.rf[6][23] ;
 wire \rvsingle.dp.rf.rf[6][24] ;
 wire \rvsingle.dp.rf.rf[6][25] ;
 wire \rvsingle.dp.rf.rf[6][26] ;
 wire \rvsingle.dp.rf.rf[6][27] ;
 wire \rvsingle.dp.rf.rf[6][28] ;
 wire \rvsingle.dp.rf.rf[6][29] ;
 wire \rvsingle.dp.rf.rf[6][2] ;
 wire \rvsingle.dp.rf.rf[6][30] ;
 wire \rvsingle.dp.rf.rf[6][31] ;
 wire \rvsingle.dp.rf.rf[6][3] ;
 wire \rvsingle.dp.rf.rf[6][4] ;
 wire \rvsingle.dp.rf.rf[6][5] ;
 wire \rvsingle.dp.rf.rf[6][6] ;
 wire \rvsingle.dp.rf.rf[6][7] ;
 wire \rvsingle.dp.rf.rf[6][8] ;
 wire \rvsingle.dp.rf.rf[6][9] ;
 wire \rvsingle.dp.rf.rf[7][0] ;
 wire \rvsingle.dp.rf.rf[7][10] ;
 wire \rvsingle.dp.rf.rf[7][11] ;
 wire \rvsingle.dp.rf.rf[7][12] ;
 wire \rvsingle.dp.rf.rf[7][13] ;
 wire \rvsingle.dp.rf.rf[7][14] ;
 wire \rvsingle.dp.rf.rf[7][15] ;
 wire \rvsingle.dp.rf.rf[7][16] ;
 wire \rvsingle.dp.rf.rf[7][17] ;
 wire \rvsingle.dp.rf.rf[7][18] ;
 wire \rvsingle.dp.rf.rf[7][19] ;
 wire \rvsingle.dp.rf.rf[7][1] ;
 wire \rvsingle.dp.rf.rf[7][20] ;
 wire \rvsingle.dp.rf.rf[7][21] ;
 wire \rvsingle.dp.rf.rf[7][22] ;
 wire \rvsingle.dp.rf.rf[7][23] ;
 wire \rvsingle.dp.rf.rf[7][24] ;
 wire \rvsingle.dp.rf.rf[7][25] ;
 wire \rvsingle.dp.rf.rf[7][26] ;
 wire \rvsingle.dp.rf.rf[7][27] ;
 wire \rvsingle.dp.rf.rf[7][28] ;
 wire \rvsingle.dp.rf.rf[7][29] ;
 wire \rvsingle.dp.rf.rf[7][2] ;
 wire \rvsingle.dp.rf.rf[7][30] ;
 wire \rvsingle.dp.rf.rf[7][31] ;
 wire \rvsingle.dp.rf.rf[7][3] ;
 wire \rvsingle.dp.rf.rf[7][4] ;
 wire \rvsingle.dp.rf.rf[7][5] ;
 wire \rvsingle.dp.rf.rf[7][6] ;
 wire \rvsingle.dp.rf.rf[7][7] ;
 wire \rvsingle.dp.rf.rf[7][8] ;
 wire \rvsingle.dp.rf.rf[7][9] ;
 wire \rvsingle.dp.rf.rf[8][0] ;
 wire \rvsingle.dp.rf.rf[8][10] ;
 wire \rvsingle.dp.rf.rf[8][11] ;
 wire \rvsingle.dp.rf.rf[8][12] ;
 wire \rvsingle.dp.rf.rf[8][13] ;
 wire \rvsingle.dp.rf.rf[8][14] ;
 wire \rvsingle.dp.rf.rf[8][15] ;
 wire \rvsingle.dp.rf.rf[8][16] ;
 wire \rvsingle.dp.rf.rf[8][17] ;
 wire \rvsingle.dp.rf.rf[8][18] ;
 wire \rvsingle.dp.rf.rf[8][19] ;
 wire \rvsingle.dp.rf.rf[8][1] ;
 wire \rvsingle.dp.rf.rf[8][20] ;
 wire \rvsingle.dp.rf.rf[8][21] ;
 wire \rvsingle.dp.rf.rf[8][22] ;
 wire \rvsingle.dp.rf.rf[8][23] ;
 wire \rvsingle.dp.rf.rf[8][24] ;
 wire \rvsingle.dp.rf.rf[8][25] ;
 wire \rvsingle.dp.rf.rf[8][26] ;
 wire \rvsingle.dp.rf.rf[8][27] ;
 wire \rvsingle.dp.rf.rf[8][28] ;
 wire \rvsingle.dp.rf.rf[8][29] ;
 wire \rvsingle.dp.rf.rf[8][2] ;
 wire \rvsingle.dp.rf.rf[8][30] ;
 wire \rvsingle.dp.rf.rf[8][31] ;
 wire \rvsingle.dp.rf.rf[8][3] ;
 wire \rvsingle.dp.rf.rf[8][4] ;
 wire \rvsingle.dp.rf.rf[8][5] ;
 wire \rvsingle.dp.rf.rf[8][6] ;
 wire \rvsingle.dp.rf.rf[8][7] ;
 wire \rvsingle.dp.rf.rf[8][8] ;
 wire \rvsingle.dp.rf.rf[8][9] ;
 wire \rvsingle.dp.rf.rf[9][0] ;
 wire \rvsingle.dp.rf.rf[9][10] ;
 wire \rvsingle.dp.rf.rf[9][11] ;
 wire \rvsingle.dp.rf.rf[9][12] ;
 wire \rvsingle.dp.rf.rf[9][13] ;
 wire \rvsingle.dp.rf.rf[9][14] ;
 wire \rvsingle.dp.rf.rf[9][15] ;
 wire \rvsingle.dp.rf.rf[9][16] ;
 wire \rvsingle.dp.rf.rf[9][17] ;
 wire \rvsingle.dp.rf.rf[9][18] ;
 wire \rvsingle.dp.rf.rf[9][19] ;
 wire \rvsingle.dp.rf.rf[9][1] ;
 wire \rvsingle.dp.rf.rf[9][20] ;
 wire \rvsingle.dp.rf.rf[9][21] ;
 wire \rvsingle.dp.rf.rf[9][22] ;
 wire \rvsingle.dp.rf.rf[9][23] ;
 wire \rvsingle.dp.rf.rf[9][24] ;
 wire \rvsingle.dp.rf.rf[9][25] ;
 wire \rvsingle.dp.rf.rf[9][26] ;
 wire \rvsingle.dp.rf.rf[9][27] ;
 wire \rvsingle.dp.rf.rf[9][28] ;
 wire \rvsingle.dp.rf.rf[9][29] ;
 wire \rvsingle.dp.rf.rf[9][2] ;
 wire \rvsingle.dp.rf.rf[9][30] ;
 wire \rvsingle.dp.rf.rf[9][31] ;
 wire \rvsingle.dp.rf.rf[9][3] ;
 wire \rvsingle.dp.rf.rf[9][4] ;
 wire \rvsingle.dp.rf.rf[9][5] ;
 wire \rvsingle.dp.rf.rf[9][6] ;
 wire \rvsingle.dp.rf.rf[9][7] ;
 wire \rvsingle.dp.rf.rf[9][8] ;
 wire \rvsingle.dp.rf.rf[9][9] ;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;

 sky130_fd_sc_hd__inv_2 _06134_ (.A(PC[1]),
    .Y(_01058_));
 sky130_fd_sc_hd__nand2_2 _06135_ (.A(Instr[13]),
    .B(Instr[14]),
    .Y(_01059_));
 sky130_fd_sc_hd__and2b_2 _06136_ (.A_N(Instr[12]),
    .B(Instr[13]),
    .X(_01060_));
 sky130_fd_sc_hd__and2b_2 _06137_ (.A_N(Instr[6]),
    .B(Instr[4]),
    .X(_01061_));
 sky130_fd_sc_hd__nor2_2 _06138_ (.A(Instr[3]),
    .B(Instr[2]),
    .Y(_01062_));
 sky130_fd_sc_hd__nand4_2 _06139_ (.A(Instr[1]),
    .B(Instr[0]),
    .C(_01061_),
    .D(_01062_),
    .Y(_01063_));
 sky130_fd_sc_hd__a311oi_2 _06140_ (.A1(Instr[30]),
    .A2(Instr[5]),
    .A3(_01059_),
    .B1(_01060_),
    .C1(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__buf_1 _06141_ (.A(_01064_),
    .X(_01065_));
 sky130_fd_sc_hd__buf_1 _06142_ (.A(_01065_),
    .X(_01066_));
 sky130_fd_sc_hd__buf_1 _06143_ (.A(Instr[6]),
    .X(_01067_));
 sky130_fd_sc_hd__nand4b_2 _06144_ (.A_N(Instr[4]),
    .B(Instr[1]),
    .C(Instr[0]),
    .D(Instr[5]),
    .Y(_01068_));
 sky130_fd_sc_hd__nor3_2 _06145_ (.A(Instr[3]),
    .B(Instr[2]),
    .C(_01068_),
    .Y(_01069_));
 sky130_fd_sc_hd__and2_2 _06146_ (.A(Instr[1]),
    .B(Instr[0]),
    .X(_01070_));
 sky130_fd_sc_hd__buf_1 _06147_ (.A(_01070_),
    .X(_01071_));
 sky130_fd_sc_hd__and3_2 _06148_ (.A(_01071_),
    .B(_01061_),
    .C(_01062_),
    .X(_01072_));
 sky130_fd_sc_hd__a21oi_2 _06149_ (.A1(_01067_),
    .A2(_01069_),
    .B1(_01072_),
    .Y(_01073_));
 sky130_fd_sc_hd__buf_1 _06150_ (.A(_01073_),
    .X(_01074_));
 sky130_fd_sc_hd__buf_1 _06151_ (.A(_01074_),
    .X(_01075_));
 sky130_fd_sc_hd__nor2b_2 _06152_ (.A(Instr[4]),
    .B_N(Instr[5]),
    .Y(_01076_));
 sky130_fd_sc_hd__nand3_2 _06153_ (.A(_01076_),
    .B(_01071_),
    .C(_01062_),
    .Y(_01077_));
 sky130_fd_sc_hd__buf_1 _06154_ (.A(_01077_),
    .X(_01078_));
 sky130_fd_sc_hd__and3_2 _06155_ (.A(Instr[6]),
    .B(Instr[3]),
    .C(Instr[2]),
    .X(_01079_));
 sky130_fd_sc_hd__nand4_2 _06156_ (.A(Instr[1]),
    .B(Instr[0]),
    .C(_01076_),
    .D(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand3_2 _06157_ (.A(_01080_),
    .B(_01063_),
    .C(_01077_),
    .Y(_01081_));
 sky130_fd_sc_hd__o221a_2 _06158_ (.A1(Instr[5]),
    .A2(_01063_),
    .B1(_01078_),
    .B2(_01067_),
    .C1(_01081_),
    .X(_01082_));
 sky130_fd_sc_hd__buf_1 _06159_ (.A(_01082_),
    .X(_01083_));
 sky130_fd_sc_hd__buf_1 _06160_ (.A(_01083_),
    .X(_01084_));
 sky130_fd_sc_hd__buf_1 _06161_ (.A(_01084_),
    .X(_01085_));
 sky130_fd_sc_hd__inv_2 _06162_ (.A(Instr[20]),
    .Y(_01086_));
 sky130_fd_sc_hd__buf_1 _06163_ (.A(_01086_),
    .X(_01087_));
 sky130_fd_sc_hd__buf_1 _06164_ (.A(_01087_),
    .X(_01088_));
 sky130_fd_sc_hd__buf_1 _06165_ (.A(_01088_),
    .X(_01089_));
 sky130_fd_sc_hd__buf_1 _06166_ (.A(_01089_),
    .X(_01090_));
 sky130_fd_sc_hd__inv_2 _06167_ (.A(Instr[21]),
    .Y(_01091_));
 sky130_fd_sc_hd__buf_1 _06168_ (.A(_01091_),
    .X(_01092_));
 sky130_fd_sc_hd__buf_1 _06169_ (.A(_01092_),
    .X(_01093_));
 sky130_fd_sc_hd__buf_1 _06170_ (.A(_01093_),
    .X(_01094_));
 sky130_fd_sc_hd__buf_1 _06171_ (.A(Instr[20]),
    .X(_01095_));
 sky130_fd_sc_hd__buf_1 _06172_ (.A(_01095_),
    .X(_01096_));
 sky130_fd_sc_hd__clkbuf_2 _06173_ (.A(_01096_),
    .X(_01097_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06174_ (.A(_01097_),
    .X(_01098_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06175_ (.A(_01098_),
    .X(_01099_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06176_ (.A(_01099_),
    .X(_01100_));
 sky130_fd_sc_hd__or2_2 _06177_ (.A(_01100_),
    .B(\rvsingle.dp.rf.rf[4][30] ),
    .X(_01101_));
 sky130_fd_sc_hd__o211ai_2 _06178_ (.A1(\rvsingle.dp.rf.rf[5][30] ),
    .A2(_01090_),
    .B1(_01094_),
    .C1(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__buf_1 _06179_ (.A(Instr[21]),
    .X(_01103_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06180_ (.A(_01103_),
    .X(_01104_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06181_ (.A(_01104_),
    .X(_01105_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06182_ (.A(_01105_),
    .X(_01106_));
 sky130_fd_sc_hd__buf_1 _06183_ (.A(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__o21a_2 _06184_ (.A1(_01100_),
    .A2(\rvsingle.dp.rf.rf[6][30] ),
    .B1(_01107_),
    .X(_01108_));
 sky130_fd_sc_hd__o21ai_2 _06185_ (.A1(\rvsingle.dp.rf.rf[7][30] ),
    .A2(_01090_),
    .B1(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__buf_1 _06186_ (.A(Instr[22]),
    .X(_01110_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06187_ (.A(_01110_),
    .X(_01111_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06188_ (.A(_01111_),
    .X(_01112_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06189_ (.A(_01112_),
    .X(_01113_));
 sky130_fd_sc_hd__buf_1 _06190_ (.A(_01113_),
    .X(_01114_));
 sky130_fd_sc_hd__buf_1 _06191_ (.A(Instr[23]),
    .X(_01115_));
 sky130_fd_sc_hd__buf_1 _06192_ (.A(_01115_),
    .X(_01116_));
 sky130_fd_sc_hd__buf_1 _06193_ (.A(_01116_),
    .X(_01117_));
 sky130_fd_sc_hd__buf_1 _06194_ (.A(_01117_),
    .X(_01118_));
 sky130_fd_sc_hd__a31o_2 _06195_ (.A1(_01102_),
    .A2(_01109_),
    .A3(_01114_),
    .B1(_01118_),
    .X(_01119_));
 sky130_fd_sc_hd__buf_1 _06196_ (.A(_01107_),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_2 _06197_ (.A0(\rvsingle.dp.rf.rf[0][30] ),
    .A1(\rvsingle.dp.rf.rf[1][30] ),
    .A2(\rvsingle.dp.rf.rf[2][30] ),
    .A3(\rvsingle.dp.rf.rf[3][30] ),
    .S0(_01100_),
    .S1(_01120_),
    .X(_01121_));
 sky130_fd_sc_hd__nor2_2 _06198_ (.A(_01114_),
    .B(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__mux4_2 _06199_ (.A0(\rvsingle.dp.rf.rf[8][30] ),
    .A1(\rvsingle.dp.rf.rf[9][30] ),
    .A2(\rvsingle.dp.rf.rf[10][30] ),
    .A3(\rvsingle.dp.rf.rf[11][30] ),
    .S0(_01100_),
    .S1(_01120_),
    .X(_01123_));
 sky130_fd_sc_hd__buf_1 _06200_ (.A(Instr[20]),
    .X(_01124_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06201_ (.A(_01124_),
    .X(_01125_));
 sky130_fd_sc_hd__clkbuf_2 _06202_ (.A(_01125_),
    .X(_01126_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06203_ (.A(_01126_),
    .X(_01127_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06204_ (.A(_01127_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_2 _06205_ (.A0(\rvsingle.dp.rf.rf[12][30] ),
    .A1(\rvsingle.dp.rf.rf[13][30] ),
    .S(_01128_),
    .X(_01129_));
 sky130_fd_sc_hd__inv_2 _06206_ (.A(Instr[22]),
    .Y(_01130_));
 sky130_fd_sc_hd__buf_1 _06207_ (.A(_01130_),
    .X(_01131_));
 sky130_fd_sc_hd__buf_1 _06208_ (.A(_01131_),
    .X(_01132_));
 sky130_fd_sc_hd__buf_1 _06209_ (.A(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__buf_1 _06210_ (.A(_01133_),
    .X(_01134_));
 sky130_fd_sc_hd__buf_1 _06211_ (.A(Instr[20]),
    .X(_01135_));
 sky130_fd_sc_hd__buf_1 _06212_ (.A(_01135_),
    .X(_01136_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06213_ (.A(_01136_),
    .X(_01137_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06214_ (.A(_01137_),
    .X(_01138_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06215_ (.A(_01138_),
    .X(_01139_));
 sky130_fd_sc_hd__or2_2 _06216_ (.A(_01139_),
    .B(\rvsingle.dp.rf.rf[14][30] ),
    .X(_01140_));
 sky130_fd_sc_hd__o211a_2 _06217_ (.A1(_01090_),
    .A2(\rvsingle.dp.rf.rf[15][30] ),
    .B1(_01107_),
    .C1(_01140_),
    .X(_01141_));
 sky130_fd_sc_hd__a211o_2 _06218_ (.A1(_01129_),
    .A2(_01094_),
    .B1(_01134_),
    .C1(_01141_),
    .X(_01142_));
 sky130_fd_sc_hd__o211ai_2 _06219_ (.A1(_01114_),
    .A2(_01123_),
    .B1(_01142_),
    .C1(_01118_),
    .Y(_01143_));
 sky130_fd_sc_hd__o21ai_2 _06220_ (.A1(_01119_),
    .A2(_01122_),
    .B1(_01143_),
    .Y(_01144_));
 sky130_fd_sc_hd__buf_1 _06221_ (.A(Instr[24]),
    .X(_01145_));
 sky130_fd_sc_hd__buf_1 _06222_ (.A(_01145_),
    .X(_01146_));
 sky130_fd_sc_hd__buf_1 _06223_ (.A(_01146_),
    .X(_01147_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06224_ (.A(_01096_),
    .X(_01148_));
 sky130_fd_sc_hd__or4_2 _06225_ (.A(_01145_),
    .B(Instr[21]),
    .C(Instr[22]),
    .D(_01115_),
    .X(_01149_));
 sky130_fd_sc_hd__buf_1 _06226_ (.A(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__or2_2 _06227_ (.A(_01148_),
    .B(_01150_),
    .X(_01151_));
 sky130_fd_sc_hd__buf_1 _06228_ (.A(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__buf_1 _06229_ (.A(_01152_),
    .X(_01153_));
 sky130_fd_sc_hd__buf_1 _06230_ (.A(_01153_),
    .X(_01154_));
 sky130_fd_sc_hd__inv_2 _06231_ (.A(_01115_),
    .Y(_01155_));
 sky130_fd_sc_hd__buf_1 _06232_ (.A(_01155_),
    .X(_01156_));
 sky130_fd_sc_hd__buf_1 _06233_ (.A(_01156_),
    .X(_01157_));
 sky130_fd_sc_hd__mux4_2 _06234_ (.A0(\rvsingle.dp.rf.rf[16][30] ),
    .A1(\rvsingle.dp.rf.rf[17][30] ),
    .A2(\rvsingle.dp.rf.rf[18][30] ),
    .A3(\rvsingle.dp.rf.rf[19][30] ),
    .S0(_01128_),
    .S1(_01107_),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_2 _06235_ (.A0(\rvsingle.dp.rf.rf[20][30] ),
    .A1(\rvsingle.dp.rf.rf[21][30] ),
    .A2(\rvsingle.dp.rf.rf[22][30] ),
    .A3(\rvsingle.dp.rf.rf[23][30] ),
    .S0(_01128_),
    .S1(_01107_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_2 _06236_ (.A0(_01158_),
    .A1(_01159_),
    .S(_01114_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_2 _06237_ (.A0(\rvsingle.dp.rf.rf[28][30] ),
    .A1(\rvsingle.dp.rf.rf[29][30] ),
    .S(_01128_),
    .X(_01161_));
 sky130_fd_sc_hd__or2_2 _06238_ (.A(_01139_),
    .B(\rvsingle.dp.rf.rf[30][30] ),
    .X(_01162_));
 sky130_fd_sc_hd__o211a_2 _06239_ (.A1(_01090_),
    .A2(\rvsingle.dp.rf.rf[31][30] ),
    .B1(_01107_),
    .C1(_01162_),
    .X(_01163_));
 sky130_fd_sc_hd__a211oi_2 _06240_ (.A1(_01161_),
    .A2(_01094_),
    .B1(_01134_),
    .C1(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__mux4_2 _06241_ (.A0(\rvsingle.dp.rf.rf[24][30] ),
    .A1(\rvsingle.dp.rf.rf[25][30] ),
    .A2(\rvsingle.dp.rf.rf[26][30] ),
    .A3(\rvsingle.dp.rf.rf[27][30] ),
    .S0(_01128_),
    .S1(_01107_),
    .X(_01165_));
 sky130_fd_sc_hd__o21ai_2 _06242_ (.A1(_01114_),
    .A2(_01165_),
    .B1(_01118_),
    .Y(_01166_));
 sky130_fd_sc_hd__o21ai_2 _06243_ (.A1(_01164_),
    .A2(_01166_),
    .B1(_01147_),
    .Y(_01167_));
 sky130_fd_sc_hd__a21o_2 _06244_ (.A1(_01157_),
    .A2(_01160_),
    .B1(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__o211a_2 _06245_ (.A1(_01144_),
    .A2(_01147_),
    .B1(_01154_),
    .C1(_01168_),
    .X(WriteData[30]));
 sky130_fd_sc_hd__inv_2 _06246_ (.A(Instr[5]),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_2 _06247_ (.A(_01071_),
    .B(_01079_),
    .Y(_01170_));
 sky130_fd_sc_hd__o31a_2 _06248_ (.A1(_01169_),
    .A2(Instr[4]),
    .A3(_01170_),
    .B1(Instr[31]),
    .X(_01171_));
 sky130_fd_sc_hd__buf_1 _06249_ (.A(Instr[17]),
    .X(_01172_));
 sky130_fd_sc_hd__nand2_2 _06250_ (.A(Instr[1]),
    .B(Instr[0]),
    .Y(_01173_));
 sky130_fd_sc_hd__nand3_2 _06251_ (.A(Instr[6]),
    .B(Instr[3]),
    .C(Instr[2]),
    .Y(_01174_));
 sky130_fd_sc_hd__nor2_2 _06252_ (.A(_01173_),
    .B(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__and3_2 _06253_ (.A(_01172_),
    .B(_01076_),
    .C(_01175_),
    .X(_01176_));
 sky130_fd_sc_hd__o221ai_2 _06254_ (.A1(Instr[5]),
    .A2(_01063_),
    .B1(_01078_),
    .B2(_01067_),
    .C1(_01081_),
    .Y(_01177_));
 sky130_fd_sc_hd__buf_1 _06255_ (.A(_01177_),
    .X(_01178_));
 sky130_fd_sc_hd__o21a_2 _06256_ (.A1(_01171_),
    .A2(_01176_),
    .B1(_01178_),
    .X(_01179_));
 sky130_fd_sc_hd__buf_1 _06257_ (.A(_01179_),
    .X(_01180_));
 sky130_fd_sc_hd__a21o_2 _06258_ (.A1(_01085_),
    .A2(WriteData[30]),
    .B1(_01180_),
    .X(_01181_));
 sky130_fd_sc_hd__or3b_2 _06259_ (.A(_01066_),
    .B(_01075_),
    .C_N(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__nor2_2 _06260_ (.A(_01064_),
    .B(_01073_),
    .Y(_01183_));
 sky130_fd_sc_hd__buf_1 _06261_ (.A(_01183_),
    .X(_01184_));
 sky130_fd_sc_hd__buf_1 _06262_ (.A(_01184_),
    .X(_01185_));
 sky130_fd_sc_hd__a211o_2 _06263_ (.A1(_01085_),
    .A2(WriteData[30]),
    .B1(_01180_),
    .C1(_01185_),
    .X(_01186_));
 sky130_fd_sc_hd__buf_1 _06264_ (.A(Instr[19]),
    .X(_01187_));
 sky130_fd_sc_hd__buf_1 _06265_ (.A(_01187_),
    .X(_01188_));
 sky130_fd_sc_hd__buf_1 _06266_ (.A(_01188_),
    .X(_01189_));
 sky130_fd_sc_hd__buf_1 _06267_ (.A(Instr[15]),
    .X(_01190_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06268_ (.A(_01190_),
    .X(_01191_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06269_ (.A(_01191_),
    .X(_01192_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06270_ (.A(_01192_),
    .X(_01193_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06271_ (.A(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__buf_1 _06272_ (.A(_01194_),
    .X(_01195_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06273_ (.A(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__buf_1 _06274_ (.A(Instr[16]),
    .X(_01197_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06275_ (.A(_01197_),
    .X(_01198_));
 sky130_fd_sc_hd__clkbuf_2 _06276_ (.A(_01198_),
    .X(_01199_));
 sky130_fd_sc_hd__clkbuf_4 _06277_ (.A(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06278_ (.A(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06279_ (.A(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06280_ (.A(_01202_),
    .X(_01203_));
 sky130_fd_sc_hd__mux4_2 _06281_ (.A0(\rvsingle.dp.rf.rf[12][30] ),
    .A1(\rvsingle.dp.rf.rf[13][30] ),
    .A2(\rvsingle.dp.rf.rf[14][30] ),
    .A3(\rvsingle.dp.rf.rf[15][30] ),
    .S0(_01196_),
    .S1(_01203_),
    .X(_01204_));
 sky130_fd_sc_hd__mux4_2 _06282_ (.A0(\rvsingle.dp.rf.rf[8][30] ),
    .A1(\rvsingle.dp.rf.rf[9][30] ),
    .A2(\rvsingle.dp.rf.rf[10][30] ),
    .A3(\rvsingle.dp.rf.rf[11][30] ),
    .S0(_01196_),
    .S1(_01203_),
    .X(_01205_));
 sky130_fd_sc_hd__inv_2 _06283_ (.A(Instr[17]),
    .Y(_01206_));
 sky130_fd_sc_hd__buf_1 _06284_ (.A(_01206_),
    .X(_01207_));
 sky130_fd_sc_hd__buf_1 _06285_ (.A(_01207_),
    .X(_01208_));
 sky130_fd_sc_hd__buf_1 _06286_ (.A(_01208_),
    .X(_01209_));
 sky130_fd_sc_hd__buf_1 _06287_ (.A(_01209_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_2 _06288_ (.A0(_01204_),
    .A1(_01205_),
    .S(_01210_),
    .X(_01211_));
 sky130_fd_sc_hd__mux4_2 _06289_ (.A0(\rvsingle.dp.rf.rf[4][30] ),
    .A1(\rvsingle.dp.rf.rf[5][30] ),
    .A2(\rvsingle.dp.rf.rf[6][30] ),
    .A3(\rvsingle.dp.rf.rf[7][30] ),
    .S0(_01196_),
    .S1(_01203_),
    .X(_01212_));
 sky130_fd_sc_hd__mux4_2 _06290_ (.A0(\rvsingle.dp.rf.rf[0][30] ),
    .A1(\rvsingle.dp.rf.rf[1][30] ),
    .A2(\rvsingle.dp.rf.rf[2][30] ),
    .A3(\rvsingle.dp.rf.rf[3][30] ),
    .S0(_01196_),
    .S1(_01203_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_2 _06291_ (.A0(_01212_),
    .A1(_01213_),
    .S(_01210_),
    .X(_01214_));
 sky130_fd_sc_hd__buf_1 _06292_ (.A(Instr[18]),
    .X(_01215_));
 sky130_fd_sc_hd__inv_2 _06293_ (.A(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__buf_1 _06294_ (.A(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__buf_1 _06295_ (.A(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__buf_1 _06296_ (.A(_01218_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_2 _06297_ (.A0(_01211_),
    .A1(_01214_),
    .S(_01219_),
    .X(_01220_));
 sky130_fd_sc_hd__buf_1 _06298_ (.A(_01215_),
    .X(_01221_));
 sky130_fd_sc_hd__buf_1 _06299_ (.A(_01221_),
    .X(_01222_));
 sky130_fd_sc_hd__buf_1 _06300_ (.A(_01222_),
    .X(_01223_));
 sky130_fd_sc_hd__buf_1 _06301_ (.A(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06302_ (.A(_01195_),
    .X(_01225_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06303_ (.A(_01203_),
    .X(_01226_));
 sky130_fd_sc_hd__mux4_2 _06304_ (.A0(\rvsingle.dp.rf.rf[20][30] ),
    .A1(\rvsingle.dp.rf.rf[21][30] ),
    .A2(\rvsingle.dp.rf.rf[22][30] ),
    .A3(\rvsingle.dp.rf.rf[23][30] ),
    .S0(_01225_),
    .S1(_01226_),
    .X(_01227_));
 sky130_fd_sc_hd__nor2_2 _06305_ (.A(_01210_),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__buf_1 _06306_ (.A(_01172_),
    .X(_01229_));
 sky130_fd_sc_hd__buf_1 _06307_ (.A(_01229_),
    .X(_01230_));
 sky130_fd_sc_hd__buf_1 _06308_ (.A(_01230_),
    .X(_01231_));
 sky130_fd_sc_hd__buf_1 _06309_ (.A(_01231_),
    .X(_01232_));
 sky130_fd_sc_hd__mux4_2 _06310_ (.A0(\rvsingle.dp.rf.rf[16][30] ),
    .A1(\rvsingle.dp.rf.rf[17][30] ),
    .A2(\rvsingle.dp.rf.rf[18][30] ),
    .A3(\rvsingle.dp.rf.rf[19][30] ),
    .S0(_01225_),
    .S1(_01226_),
    .X(_01233_));
 sky130_fd_sc_hd__nor2_2 _06311_ (.A(_01232_),
    .B(_01233_),
    .Y(_01234_));
 sky130_fd_sc_hd__mux4_2 _06312_ (.A0(\rvsingle.dp.rf.rf[24][30] ),
    .A1(\rvsingle.dp.rf.rf[25][30] ),
    .A2(\rvsingle.dp.rf.rf[26][30] ),
    .A3(\rvsingle.dp.rf.rf[27][30] ),
    .S0(_01225_),
    .S1(_01226_),
    .X(_01235_));
 sky130_fd_sc_hd__mux4_2 _06313_ (.A0(\rvsingle.dp.rf.rf[28][30] ),
    .A1(\rvsingle.dp.rf.rf[29][30] ),
    .A2(\rvsingle.dp.rf.rf[30][30] ),
    .A3(\rvsingle.dp.rf.rf[31][30] ),
    .S0(_01196_),
    .S1(_01203_),
    .X(_01236_));
 sky130_fd_sc_hd__o21a_2 _06314_ (.A1(_01210_),
    .A2(_01236_),
    .B1(_01224_),
    .X(_01237_));
 sky130_fd_sc_hd__o21ai_2 _06315_ (.A1(_01232_),
    .A2(_01235_),
    .B1(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__o311ai_2 _06316_ (.A1(_01224_),
    .A2(_01228_),
    .A3(_01234_),
    .B1(_01189_),
    .C1(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06317_ (.A(_01190_),
    .X(_01240_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06318_ (.A(_01240_),
    .X(_01241_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06319_ (.A(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06320_ (.A(_01197_),
    .X(_01243_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06321_ (.A(_01243_),
    .X(_01244_));
 sky130_fd_sc_hd__or3_2 _06322_ (.A(Instr[17]),
    .B(_01215_),
    .C(Instr[19]),
    .X(_01245_));
 sky130_fd_sc_hd__or3_2 _06323_ (.A(_01242_),
    .B(_01244_),
    .C(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06324_ (.A(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06325_ (.A(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__o211a_2 _06326_ (.A1(_01189_),
    .A2(_01220_),
    .B1(_01239_),
    .C1(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__nand3_2 _06327_ (.A(_01182_),
    .B(_01186_),
    .C(_01249_),
    .Y(_01250_));
 sky130_fd_sc_hd__or2_2 _06328_ (.A(_01099_),
    .B(\rvsingle.dp.rf.rf[0][29] ),
    .X(_01251_));
 sky130_fd_sc_hd__o211ai_2 _06329_ (.A1(\rvsingle.dp.rf.rf[1][29] ),
    .A2(_01089_),
    .B1(_01093_),
    .C1(_01251_),
    .Y(_01252_));
 sky130_fd_sc_hd__mux2_2 _06330_ (.A0(\rvsingle.dp.rf.rf[2][29] ),
    .A1(\rvsingle.dp.rf.rf[3][29] ),
    .S(_01138_),
    .X(_01253_));
 sky130_fd_sc_hd__a21oi_2 _06331_ (.A1(_01107_),
    .A2(_01253_),
    .B1(_01113_),
    .Y(_01254_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06332_ (.A(_01095_),
    .X(_01255_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06333_ (.A(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06334_ (.A(_01256_),
    .X(_01257_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06335_ (.A(Instr[21]),
    .X(_01258_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06336_ (.A(_01258_),
    .X(_01259_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06337_ (.A(_01259_),
    .X(_01260_));
 sky130_fd_sc_hd__buf_1 _06338_ (.A(_01260_),
    .X(_01261_));
 sky130_fd_sc_hd__mux4_2 _06339_ (.A0(\rvsingle.dp.rf.rf[4][29] ),
    .A1(\rvsingle.dp.rf.rf[5][29] ),
    .A2(\rvsingle.dp.rf.rf[6][29] ),
    .A3(\rvsingle.dp.rf.rf[7][29] ),
    .S0(_01257_),
    .S1(_01261_),
    .X(_01262_));
 sky130_fd_sc_hd__o2bb2a_2 _06340_ (.A1_N(_01252_),
    .A2_N(_01254_),
    .B1(_01133_),
    .B2(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__mux4_2 _06341_ (.A0(\rvsingle.dp.rf.rf[8][29] ),
    .A1(\rvsingle.dp.rf.rf[9][29] ),
    .A2(\rvsingle.dp.rf.rf[10][29] ),
    .A3(\rvsingle.dp.rf.rf[11][29] ),
    .S0(_01127_),
    .S1(_01261_),
    .X(_01264_));
 sky130_fd_sc_hd__or2_2 _06342_ (.A(_01138_),
    .B(\rvsingle.dp.rf.rf[12][29] ),
    .X(_01265_));
 sky130_fd_sc_hd__o211a_2 _06343_ (.A1(\rvsingle.dp.rf.rf[13][29] ),
    .A2(_01089_),
    .B1(_01093_),
    .C1(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__buf_1 _06344_ (.A(_01135_),
    .X(_01267_));
 sky130_fd_sc_hd__buf_1 _06345_ (.A(_01267_),
    .X(_01268_));
 sky130_fd_sc_hd__buf_1 _06346_ (.A(_01268_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_2 _06347_ (.A0(\rvsingle.dp.rf.rf[14][29] ),
    .A1(\rvsingle.dp.rf.rf[15][29] ),
    .S(_01269_),
    .X(_01270_));
 sky130_fd_sc_hd__a21o_2 _06348_ (.A1(_01261_),
    .A2(_01270_),
    .B1(_01133_),
    .X(_01271_));
 sky130_fd_sc_hd__o221a_2 _06349_ (.A1(_01113_),
    .A2(_01264_),
    .B1(_01266_),
    .B2(_01271_),
    .C1(_01118_),
    .X(_01272_));
 sky130_fd_sc_hd__a21o_2 _06350_ (.A1(_01157_),
    .A2(_01263_),
    .B1(_01272_),
    .X(_01273_));
 sky130_fd_sc_hd__mux4_2 _06351_ (.A0(\rvsingle.dp.rf.rf[16][29] ),
    .A1(\rvsingle.dp.rf.rf[17][29] ),
    .A2(\rvsingle.dp.rf.rf[18][29] ),
    .A3(\rvsingle.dp.rf.rf[19][29] ),
    .S0(_01139_),
    .S1(_01261_),
    .X(_01274_));
 sky130_fd_sc_hd__nor2_2 _06352_ (.A(_01113_),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__mux2_2 _06353_ (.A0(\rvsingle.dp.rf.rf[20][29] ),
    .A1(\rvsingle.dp.rf.rf[21][29] ),
    .S(_01139_),
    .X(_01276_));
 sky130_fd_sc_hd__or2_2 _06354_ (.A(_01099_),
    .B(\rvsingle.dp.rf.rf[22][29] ),
    .X(_01277_));
 sky130_fd_sc_hd__o211a_2 _06355_ (.A1(_01089_),
    .A2(\rvsingle.dp.rf.rf[23][29] ),
    .B1(_01107_),
    .C1(_01277_),
    .X(_01278_));
 sky130_fd_sc_hd__a211oi_2 _06356_ (.A1(_01276_),
    .A2(_01094_),
    .B1(_01134_),
    .C1(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__o21a_2 _06357_ (.A1(_01139_),
    .A2(\rvsingle.dp.rf.rf[26][29] ),
    .B1(_01261_),
    .X(_01280_));
 sky130_fd_sc_hd__o21ai_2 _06358_ (.A1(\rvsingle.dp.rf.rf[27][29] ),
    .A2(_01090_),
    .B1(_01280_),
    .Y(_01281_));
 sky130_fd_sc_hd__or2_2 _06359_ (.A(_01099_),
    .B(\rvsingle.dp.rf.rf[24][29] ),
    .X(_01282_));
 sky130_fd_sc_hd__o211ai_2 _06360_ (.A1(\rvsingle.dp.rf.rf[25][29] ),
    .A2(_01090_),
    .B1(_01094_),
    .C1(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hd__mux4_2 _06361_ (.A0(\rvsingle.dp.rf.rf[28][29] ),
    .A1(\rvsingle.dp.rf.rf[29][29] ),
    .A2(\rvsingle.dp.rf.rf[30][29] ),
    .A3(\rvsingle.dp.rf.rf[31][29] ),
    .S0(_01138_),
    .S1(_01106_),
    .X(_01284_));
 sky130_fd_sc_hd__o21ai_2 _06362_ (.A1(_01133_),
    .A2(_01284_),
    .B1(_01117_),
    .Y(_01285_));
 sky130_fd_sc_hd__a31o_2 _06363_ (.A1(_01134_),
    .A2(_01281_),
    .A3(_01283_),
    .B1(_01285_),
    .X(_01286_));
 sky130_fd_sc_hd__o311ai_2 _06364_ (.A1(_01118_),
    .A2(_01275_),
    .A3(_01279_),
    .B1(_01286_),
    .C1(_01147_),
    .Y(_01287_));
 sky130_fd_sc_hd__o211a_2 _06365_ (.A1(_01147_),
    .A2(_01273_),
    .B1(_01287_),
    .C1(_01154_),
    .X(WriteData[29]));
 sky130_fd_sc_hd__a211o_2 _06366_ (.A1(_01085_),
    .A2(WriteData[29]),
    .B1(_01180_),
    .C1(_01184_),
    .X(_01288_));
 sky130_fd_sc_hd__a21o_2 _06367_ (.A1(_01085_),
    .A2(WriteData[29]),
    .B1(_01180_),
    .X(_01289_));
 sky130_fd_sc_hd__nand2_2 _06368_ (.A(_01289_),
    .B(_01184_),
    .Y(_01290_));
 sky130_fd_sc_hd__mux4_2 _06369_ (.A0(\rvsingle.dp.rf.rf[4][29] ),
    .A1(\rvsingle.dp.rf.rf[5][29] ),
    .A2(\rvsingle.dp.rf.rf[6][29] ),
    .A3(\rvsingle.dp.rf.rf[7][29] ),
    .S0(_01195_),
    .S1(_01202_),
    .X(_01291_));
 sky130_fd_sc_hd__nor2_2 _06370_ (.A(_01210_),
    .B(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hd__inv_2 _06371_ (.A(Instr[15]),
    .Y(_01293_));
 sky130_fd_sc_hd__buf_1 _06372_ (.A(_01293_),
    .X(_01294_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06373_ (.A(_01294_),
    .X(_01295_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06374_ (.A(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__buf_1 _06375_ (.A(_01296_),
    .X(_01297_));
 sky130_fd_sc_hd__buf_1 _06376_ (.A(_01297_),
    .X(_01298_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06377_ (.A(_01197_),
    .X(_01299_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06378_ (.A(_01299_),
    .X(_01300_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06379_ (.A(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06380_ (.A(_01301_),
    .X(_01302_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06381_ (.A(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__o21a_2 _06382_ (.A1(_01195_),
    .A2(\rvsingle.dp.rf.rf[2][29] ),
    .B1(_01303_),
    .X(_01304_));
 sky130_fd_sc_hd__o21ai_2 _06383_ (.A1(\rvsingle.dp.rf.rf[3][29] ),
    .A2(_01298_),
    .B1(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__inv_2 _06384_ (.A(Instr[16]),
    .Y(_01306_));
 sky130_fd_sc_hd__buf_1 _06385_ (.A(_01306_),
    .X(_01307_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06386_ (.A(_01307_),
    .X(_01308_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06387_ (.A(_01308_),
    .X(_01309_));
 sky130_fd_sc_hd__buf_1 _06388_ (.A(_01309_),
    .X(_01310_));
 sky130_fd_sc_hd__buf_1 _06389_ (.A(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__or2_2 _06390_ (.A(_01195_),
    .B(\rvsingle.dp.rf.rf[0][29] ),
    .X(_01312_));
 sky130_fd_sc_hd__o211ai_2 _06391_ (.A1(\rvsingle.dp.rf.rf[1][29] ),
    .A2(_01298_),
    .B1(_01311_),
    .C1(_01312_),
    .Y(_01313_));
 sky130_fd_sc_hd__and3_2 _06392_ (.A(_01210_),
    .B(_01305_),
    .C(_01313_),
    .X(_01314_));
 sky130_fd_sc_hd__inv_2 _06393_ (.A(Instr[19]),
    .Y(_01315_));
 sky130_fd_sc_hd__buf_1 _06394_ (.A(_01315_),
    .X(_01316_));
 sky130_fd_sc_hd__buf_1 _06395_ (.A(_01316_),
    .X(_01317_));
 sky130_fd_sc_hd__mux4_2 _06396_ (.A0(\rvsingle.dp.rf.rf[8][29] ),
    .A1(\rvsingle.dp.rf.rf[9][29] ),
    .A2(\rvsingle.dp.rf.rf[10][29] ),
    .A3(\rvsingle.dp.rf.rf[11][29] ),
    .S0(_01195_),
    .S1(_01202_),
    .X(_01318_));
 sky130_fd_sc_hd__or2_2 _06397_ (.A(_01195_),
    .B(\rvsingle.dp.rf.rf[12][29] ),
    .X(_01319_));
 sky130_fd_sc_hd__o211a_2 _06398_ (.A1(\rvsingle.dp.rf.rf[13][29] ),
    .A2(_01298_),
    .B1(_01311_),
    .C1(_01319_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_2 _06399_ (.A0(\rvsingle.dp.rf.rf[14][29] ),
    .A1(\rvsingle.dp.rf.rf[15][29] ),
    .S(_01195_),
    .X(_01321_));
 sky130_fd_sc_hd__a21o_2 _06400_ (.A1(_01202_),
    .A2(_01321_),
    .B1(_01209_),
    .X(_01322_));
 sky130_fd_sc_hd__o221ai_2 _06401_ (.A1(_01232_),
    .A2(_01318_),
    .B1(_01320_),
    .B2(_01322_),
    .C1(_01224_),
    .Y(_01323_));
 sky130_fd_sc_hd__o311ai_2 _06402_ (.A1(_01224_),
    .A2(_01292_),
    .A3(_01314_),
    .B1(_01317_),
    .C1(_01323_),
    .Y(_01324_));
 sky130_fd_sc_hd__mux4_2 _06403_ (.A0(\rvsingle.dp.rf.rf[24][29] ),
    .A1(\rvsingle.dp.rf.rf[25][29] ),
    .A2(\rvsingle.dp.rf.rf[26][29] ),
    .A3(\rvsingle.dp.rf.rf[27][29] ),
    .S0(_01194_),
    .S1(_01303_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_2 _06404_ (.A0(\rvsingle.dp.rf.rf[28][29] ),
    .A1(\rvsingle.dp.rf.rf[29][29] ),
    .S(_01194_),
    .X(_01326_));
 sky130_fd_sc_hd__buf_1 _06405_ (.A(Instr[15]),
    .X(_01327_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06406_ (.A(_01327_),
    .X(_01328_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06407_ (.A(_01328_),
    .X(_01329_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06408_ (.A(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__or2_2 _06409_ (.A(_01330_),
    .B(\rvsingle.dp.rf.rf[30][29] ),
    .X(_01331_));
 sky130_fd_sc_hd__o211a_2 _06410_ (.A1(_01297_),
    .A2(\rvsingle.dp.rf.rf[31][29] ),
    .B1(_01201_),
    .C1(_01331_),
    .X(_01332_));
 sky130_fd_sc_hd__a211o_2 _06411_ (.A1(_01326_),
    .A2(_01311_),
    .B1(_01209_),
    .C1(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__o211a_2 _06412_ (.A1(_01231_),
    .A2(_01325_),
    .B1(_01333_),
    .C1(_01223_),
    .X(_01334_));
 sky130_fd_sc_hd__clkbuf_4 _06413_ (.A(_01240_),
    .X(_01335_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06414_ (.A(_01335_),
    .X(_01336_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06415_ (.A(_01336_),
    .X(_01337_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06416_ (.A(_01337_),
    .X(_01338_));
 sky130_fd_sc_hd__mux4_2 _06417_ (.A0(\rvsingle.dp.rf.rf[16][29] ),
    .A1(\rvsingle.dp.rf.rf[17][29] ),
    .A2(\rvsingle.dp.rf.rf[18][29] ),
    .A3(\rvsingle.dp.rf.rf[19][29] ),
    .S0(_01338_),
    .S1(_01303_),
    .X(_01339_));
 sky130_fd_sc_hd__or2_2 _06418_ (.A(_01337_),
    .B(\rvsingle.dp.rf.rf[20][29] ),
    .X(_01340_));
 sky130_fd_sc_hd__o211ai_2 _06419_ (.A1(\rvsingle.dp.rf.rf[21][29] ),
    .A2(_01297_),
    .B1(_01310_),
    .C1(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__o21a_2 _06420_ (.A1(_01337_),
    .A2(\rvsingle.dp.rf.rf[22][29] ),
    .B1(_01302_),
    .X(_01342_));
 sky130_fd_sc_hd__o21ai_2 _06421_ (.A1(\rvsingle.dp.rf.rf[23][29] ),
    .A2(_01297_),
    .B1(_01342_),
    .Y(_01343_));
 sky130_fd_sc_hd__a31o_2 _06422_ (.A1(_01341_),
    .A2(_01231_),
    .A3(_01343_),
    .B1(_01222_),
    .X(_01344_));
 sky130_fd_sc_hd__o21ba_2 _06423_ (.A1(_01231_),
    .A2(_01339_),
    .B1_N(_01344_),
    .X(_01345_));
 sky130_fd_sc_hd__or3_2 _06424_ (.A(_01317_),
    .B(_01334_),
    .C(_01345_),
    .X(_01346_));
 sky130_fd_sc_hd__and3_2 _06425_ (.A(_01248_),
    .B(_01324_),
    .C(_01346_),
    .X(_01347_));
 sky130_fd_sc_hd__a21oi_2 _06426_ (.A1(_01288_),
    .A2(_01290_),
    .B1(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__buf_1 _06427_ (.A(_01190_),
    .X(_01349_));
 sky130_fd_sc_hd__or4_2 _06428_ (.A(_01349_),
    .B(Instr[17]),
    .C(_01215_),
    .D(Instr[19]),
    .X(_01350_));
 sky130_fd_sc_hd__buf_1 _06429_ (.A(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__mux4_2 _06430_ (.A0(\rvsingle.dp.rf.rf[16][28] ),
    .A1(\rvsingle.dp.rf.rf[17][28] ),
    .A2(\rvsingle.dp.rf.rf[18][28] ),
    .A3(\rvsingle.dp.rf.rf[19][28] ),
    .S0(_01338_),
    .S1(_01303_),
    .X(_01352_));
 sky130_fd_sc_hd__mux4_2 _06431_ (.A0(\rvsingle.dp.rf.rf[20][28] ),
    .A1(\rvsingle.dp.rf.rf[21][28] ),
    .A2(\rvsingle.dp.rf.rf[22][28] ),
    .A3(\rvsingle.dp.rf.rf[23][28] ),
    .S0(_01338_),
    .S1(_01303_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_2 _06432_ (.A0(_01352_),
    .A1(_01353_),
    .S(_01231_),
    .X(_01354_));
 sky130_fd_sc_hd__mux4_2 _06433_ (.A0(\rvsingle.dp.rf.rf[24][28] ),
    .A1(\rvsingle.dp.rf.rf[25][28] ),
    .A2(\rvsingle.dp.rf.rf[26][28] ),
    .A3(\rvsingle.dp.rf.rf[27][28] ),
    .S0(_01338_),
    .S1(_01202_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_2 _06434_ (.A0(\rvsingle.dp.rf.rf[28][28] ),
    .A1(\rvsingle.dp.rf.rf[29][28] ),
    .S(_01194_),
    .X(_01356_));
 sky130_fd_sc_hd__or2_2 _06435_ (.A(_01337_),
    .B(\rvsingle.dp.rf.rf[30][28] ),
    .X(_01357_));
 sky130_fd_sc_hd__o211a_2 _06436_ (.A1(_01297_),
    .A2(\rvsingle.dp.rf.rf[31][28] ),
    .B1(_01303_),
    .C1(_01357_),
    .X(_01358_));
 sky130_fd_sc_hd__a211o_2 _06437_ (.A1(_01356_),
    .A2(_01311_),
    .B1(_01209_),
    .C1(_01358_),
    .X(_01359_));
 sky130_fd_sc_hd__o211a_2 _06438_ (.A1(_01232_),
    .A2(_01355_),
    .B1(_01359_),
    .C1(_01224_),
    .X(_01360_));
 sky130_fd_sc_hd__a211o_2 _06439_ (.A1(_01219_),
    .A2(_01354_),
    .B1(_01360_),
    .C1(_01317_),
    .X(_01361_));
 sky130_fd_sc_hd__or2_2 _06440_ (.A(_01195_),
    .B(\rvsingle.dp.rf.rf[0][28] ),
    .X(_01362_));
 sky130_fd_sc_hd__o211ai_2 _06441_ (.A1(\rvsingle.dp.rf.rf[1][28] ),
    .A2(_01298_),
    .B1(_01311_),
    .C1(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__mux2_2 _06442_ (.A0(\rvsingle.dp.rf.rf[2][28] ),
    .A1(\rvsingle.dp.rf.rf[3][28] ),
    .S(_01338_),
    .X(_01364_));
 sky130_fd_sc_hd__a21oi_2 _06443_ (.A1(_01202_),
    .A2(_01364_),
    .B1(_01231_),
    .Y(_01365_));
 sky130_fd_sc_hd__mux4_2 _06444_ (.A0(\rvsingle.dp.rf.rf[4][28] ),
    .A1(\rvsingle.dp.rf.rf[5][28] ),
    .A2(\rvsingle.dp.rf.rf[6][28] ),
    .A3(\rvsingle.dp.rf.rf[7][28] ),
    .S0(_01338_),
    .S1(_01202_),
    .X(_01366_));
 sky130_fd_sc_hd__o2bb2a_2 _06445_ (.A1_N(_01363_),
    .A2_N(_01365_),
    .B1(_01210_),
    .B2(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__mux4_2 _06446_ (.A0(\rvsingle.dp.rf.rf[8][28] ),
    .A1(\rvsingle.dp.rf.rf[9][28] ),
    .A2(\rvsingle.dp.rf.rf[10][28] ),
    .A3(\rvsingle.dp.rf.rf[11][28] ),
    .S0(_01338_),
    .S1(_01303_),
    .X(_01368_));
 sky130_fd_sc_hd__or2_2 _06447_ (.A(_01338_),
    .B(\rvsingle.dp.rf.rf[12][28] ),
    .X(_01369_));
 sky130_fd_sc_hd__o211a_2 _06448_ (.A1(\rvsingle.dp.rf.rf[13][28] ),
    .A2(_01298_),
    .B1(_01311_),
    .C1(_01369_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_2 _06449_ (.A0(\rvsingle.dp.rf.rf[14][28] ),
    .A1(\rvsingle.dp.rf.rf[15][28] ),
    .S(_01194_),
    .X(_01371_));
 sky130_fd_sc_hd__a21o_2 _06450_ (.A1(_01202_),
    .A2(_01371_),
    .B1(_01209_),
    .X(_01372_));
 sky130_fd_sc_hd__o221a_2 _06451_ (.A1(_01232_),
    .A2(_01368_),
    .B1(_01370_),
    .B2(_01372_),
    .C1(_01224_),
    .X(_01373_));
 sky130_fd_sc_hd__a211o_2 _06452_ (.A1(_01219_),
    .A2(_01367_),
    .B1(_01373_),
    .C1(_01189_),
    .X(_01374_));
 sky130_fd_sc_hd__o211ai_2 _06453_ (.A1(_01351_),
    .A2(_01226_),
    .B1(_01361_),
    .C1(_01374_),
    .Y(_01375_));
 sky130_fd_sc_hd__inv_2 _06454_ (.A(_01145_),
    .Y(_01376_));
 sky130_fd_sc_hd__buf_1 _06455_ (.A(_01376_),
    .X(_01377_));
 sky130_fd_sc_hd__buf_1 _06456_ (.A(_01377_),
    .X(_01378_));
 sky130_fd_sc_hd__mux4_2 _06457_ (.A0(\rvsingle.dp.rf.rf[24][28] ),
    .A1(\rvsingle.dp.rf.rf[25][28] ),
    .A2(\rvsingle.dp.rf.rf[26][28] ),
    .A3(\rvsingle.dp.rf.rf[27][28] ),
    .S0(_01099_),
    .S1(_01261_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_2 _06458_ (.A0(\rvsingle.dp.rf.rf[28][28] ),
    .A1(\rvsingle.dp.rf.rf[29][28] ),
    .S(_01127_),
    .X(_01380_));
 sky130_fd_sc_hd__buf_1 _06459_ (.A(_01095_),
    .X(_01381_));
 sky130_fd_sc_hd__buf_1 _06460_ (.A(_01381_),
    .X(_01382_));
 sky130_fd_sc_hd__buf_1 _06461_ (.A(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__or2_2 _06462_ (.A(_01383_),
    .B(\rvsingle.dp.rf.rf[30][28] ),
    .X(_01384_));
 sky130_fd_sc_hd__o211a_2 _06463_ (.A1(_01089_),
    .A2(\rvsingle.dp.rf.rf[31][28] ),
    .B1(_01106_),
    .C1(_01384_),
    .X(_01385_));
 sky130_fd_sc_hd__a211o_2 _06464_ (.A1(_01380_),
    .A2(_01093_),
    .B1(_01133_),
    .C1(_01385_),
    .X(_01386_));
 sky130_fd_sc_hd__o211a_2 _06465_ (.A1(_01113_),
    .A2(_01379_),
    .B1(_01386_),
    .C1(_01118_),
    .X(_01387_));
 sky130_fd_sc_hd__mux4_2 _06466_ (.A0(\rvsingle.dp.rf.rf[16][28] ),
    .A1(\rvsingle.dp.rf.rf[17][28] ),
    .A2(\rvsingle.dp.rf.rf[18][28] ),
    .A3(\rvsingle.dp.rf.rf[19][28] ),
    .S0(_01139_),
    .S1(_01107_),
    .X(_01388_));
 sky130_fd_sc_hd__mux4_2 _06467_ (.A0(\rvsingle.dp.rf.rf[20][28] ),
    .A1(\rvsingle.dp.rf.rf[21][28] ),
    .A2(\rvsingle.dp.rf.rf[22][28] ),
    .A3(\rvsingle.dp.rf.rf[23][28] ),
    .S0(_01138_),
    .S1(_01106_),
    .X(_01389_));
 sky130_fd_sc_hd__o21a_2 _06468_ (.A1(_01133_),
    .A2(_01389_),
    .B1(_01157_),
    .X(_01390_));
 sky130_fd_sc_hd__o21a_2 _06469_ (.A1(_01114_),
    .A2(_01388_),
    .B1(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__mux4_2 _06470_ (.A0(\rvsingle.dp.rf.rf[4][28] ),
    .A1(\rvsingle.dp.rf.rf[5][28] ),
    .A2(\rvsingle.dp.rf.rf[6][28] ),
    .A3(\rvsingle.dp.rf.rf[7][28] ),
    .S0(_01099_),
    .S1(_01261_),
    .X(_01392_));
 sky130_fd_sc_hd__or2_2 _06471_ (.A(_01099_),
    .B(\rvsingle.dp.rf.rf[2][28] ),
    .X(_01393_));
 sky130_fd_sc_hd__o211a_2 _06472_ (.A1(_01089_),
    .A2(\rvsingle.dp.rf.rf[3][28] ),
    .B1(_01261_),
    .C1(_01393_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_2 _06473_ (.A0(\rvsingle.dp.rf.rf[0][28] ),
    .A1(\rvsingle.dp.rf.rf[1][28] ),
    .S(_01127_),
    .X(_01395_));
 sky130_fd_sc_hd__a21o_2 _06474_ (.A1(_01395_),
    .A2(_01094_),
    .B1(_01113_),
    .X(_01396_));
 sky130_fd_sc_hd__o22ai_2 _06475_ (.A1(_01134_),
    .A2(_01392_),
    .B1(_01394_),
    .B2(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__mux4_2 _06476_ (.A0(\rvsingle.dp.rf.rf[12][28] ),
    .A1(\rvsingle.dp.rf.rf[13][28] ),
    .A2(\rvsingle.dp.rf.rf[14][28] ),
    .A3(\rvsingle.dp.rf.rf[15][28] ),
    .S0(_01099_),
    .S1(_01261_),
    .X(_01398_));
 sky130_fd_sc_hd__or2_2 _06477_ (.A(_01127_),
    .B(\rvsingle.dp.rf.rf[10][28] ),
    .X(_01399_));
 sky130_fd_sc_hd__o211a_2 _06478_ (.A1(_01089_),
    .A2(\rvsingle.dp.rf.rf[11][28] ),
    .B1(_01261_),
    .C1(_01399_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_2 _06479_ (.A0(\rvsingle.dp.rf.rf[8][28] ),
    .A1(\rvsingle.dp.rf.rf[9][28] ),
    .S(_01257_),
    .X(_01401_));
 sky130_fd_sc_hd__a21o_2 _06480_ (.A1(_01401_),
    .A2(_01093_),
    .B1(_01113_),
    .X(_01402_));
 sky130_fd_sc_hd__o221ai_2 _06481_ (.A1(_01134_),
    .A2(_01398_),
    .B1(_01400_),
    .B2(_01402_),
    .C1(_01118_),
    .Y(_01403_));
 sky130_fd_sc_hd__o211ai_2 _06482_ (.A1(_01118_),
    .A2(_01397_),
    .B1(_01403_),
    .C1(_01378_),
    .Y(_01404_));
 sky130_fd_sc_hd__o311a_2 _06483_ (.A1(_01378_),
    .A2(_01387_),
    .A3(_01391_),
    .B1(_01404_),
    .C1(_01154_),
    .X(WriteData[28]));
 sky130_fd_sc_hd__a21o_2 _06484_ (.A1(_01085_),
    .A2(WriteData[28]),
    .B1(_01180_),
    .X(_01405_));
 sky130_fd_sc_hd__or3b_2 _06485_ (.A(_01066_),
    .B(_01075_),
    .C_N(_01405_),
    .X(_01406_));
 sky130_fd_sc_hd__a211o_2 _06486_ (.A1(_01085_),
    .A2(WriteData[28]),
    .B1(_01180_),
    .C1(_01184_),
    .X(_01407_));
 sky130_fd_sc_hd__nand3b_2 _06487_ (.A_N(_01375_),
    .B(_01406_),
    .C(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__inv_2 _06488_ (.A(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hd__a31oi_2 _06489_ (.A1(_01347_),
    .A2(_01288_),
    .A3(_01290_),
    .B1(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__nand3_2 _06490_ (.A(_01375_),
    .B(_01406_),
    .C(_01407_),
    .Y(_01411_));
 sky130_fd_sc_hd__a21o_2 _06491_ (.A1(_01406_),
    .A2(_01407_),
    .B1(_01375_),
    .X(_01412_));
 sky130_fd_sc_hd__nand3_2 _06492_ (.A(_01347_),
    .B(_01288_),
    .C(_01290_),
    .Y(_01413_));
 sky130_fd_sc_hd__or2b_2 _06493_ (.A(_01348_),
    .B_N(_01413_),
    .X(_01414_));
 sky130_fd_sc_hd__a21o_2 _06494_ (.A1(_01411_),
    .A2(_01412_),
    .B1(_01414_),
    .X(_01415_));
 sky130_fd_sc_hd__buf_1 _06495_ (.A(_01327_),
    .X(_01416_));
 sky130_fd_sc_hd__buf_1 _06496_ (.A(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__mux4_2 _06497_ (.A0(\rvsingle.dp.rf.rf[24][21] ),
    .A1(\rvsingle.dp.rf.rf[25][21] ),
    .A2(\rvsingle.dp.rf.rf[26][21] ),
    .A3(\rvsingle.dp.rf.rf[27][21] ),
    .S0(_01417_),
    .S1(_01301_),
    .X(_01418_));
 sky130_fd_sc_hd__buf_1 _06498_ (.A(_01190_),
    .X(_01419_));
 sky130_fd_sc_hd__buf_1 _06499_ (.A(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_2 _06500_ (.A0(\rvsingle.dp.rf.rf[28][21] ),
    .A1(\rvsingle.dp.rf.rf[29][21] ),
    .S(_01420_),
    .X(_01421_));
 sky130_fd_sc_hd__buf_1 _06501_ (.A(_01206_),
    .X(_01422_));
 sky130_fd_sc_hd__buf_1 _06502_ (.A(_01293_),
    .X(_01423_));
 sky130_fd_sc_hd__buf_1 _06503_ (.A(_01423_),
    .X(_01424_));
 sky130_fd_sc_hd__buf_1 _06504_ (.A(Instr[15]),
    .X(_01425_));
 sky130_fd_sc_hd__buf_1 _06505_ (.A(_01425_),
    .X(_01426_));
 sky130_fd_sc_hd__buf_1 _06506_ (.A(_01197_),
    .X(_01427_));
 sky130_fd_sc_hd__o21a_2 _06507_ (.A1(_01426_),
    .A2(\rvsingle.dp.rf.rf[30][21] ),
    .B1(_01427_),
    .X(_01428_));
 sky130_fd_sc_hd__o21a_2 _06508_ (.A1(_01424_),
    .A2(\rvsingle.dp.rf.rf[31][21] ),
    .B1(_01428_),
    .X(_01429_));
 sky130_fd_sc_hd__a211o_2 _06509_ (.A1(_01421_),
    .A2(_01309_),
    .B1(_01422_),
    .C1(_01429_),
    .X(_01430_));
 sky130_fd_sc_hd__o211ai_2 _06510_ (.A1(_01230_),
    .A2(_01418_),
    .B1(_01430_),
    .C1(_01222_),
    .Y(_01431_));
 sky130_fd_sc_hd__buf_1 _06511_ (.A(_01426_),
    .X(_01432_));
 sky130_fd_sc_hd__buf_1 _06512_ (.A(_01299_),
    .X(_01433_));
 sky130_fd_sc_hd__buf_1 _06513_ (.A(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__mux4_2 _06514_ (.A0(\rvsingle.dp.rf.rf[16][21] ),
    .A1(\rvsingle.dp.rf.rf[17][21] ),
    .A2(\rvsingle.dp.rf.rf[18][21] ),
    .A3(\rvsingle.dp.rf.rf[19][21] ),
    .S0(_01432_),
    .S1(_01434_),
    .X(_01435_));
 sky130_fd_sc_hd__buf_1 _06515_ (.A(_01306_),
    .X(_01436_));
 sky130_fd_sc_hd__buf_1 _06516_ (.A(_01436_),
    .X(_01437_));
 sky130_fd_sc_hd__or2_2 _06517_ (.A(_01192_),
    .B(\rvsingle.dp.rf.rf[20][21] ),
    .X(_01438_));
 sky130_fd_sc_hd__o211ai_2 _06518_ (.A1(\rvsingle.dp.rf.rf[21][21] ),
    .A2(_01296_),
    .B1(_01437_),
    .C1(_01438_),
    .Y(_01439_));
 sky130_fd_sc_hd__buf_1 _06519_ (.A(_01294_),
    .X(_01440_));
 sky130_fd_sc_hd__buf_1 _06520_ (.A(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__or2_2 _06521_ (.A(_01420_),
    .B(\rvsingle.dp.rf.rf[22][21] ),
    .X(_01442_));
 sky130_fd_sc_hd__o211ai_2 _06522_ (.A1(_01441_),
    .A2(\rvsingle.dp.rf.rf[23][21] ),
    .B1(_01301_),
    .C1(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__buf_1 _06523_ (.A(_01172_),
    .X(_01444_));
 sky130_fd_sc_hd__buf_1 _06524_ (.A(_01444_),
    .X(_01445_));
 sky130_fd_sc_hd__buf_1 _06525_ (.A(_01215_),
    .X(_01446_));
 sky130_fd_sc_hd__buf_1 _06526_ (.A(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__a31oi_2 _06527_ (.A1(_01439_),
    .A2(_01443_),
    .A3(_01445_),
    .B1(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__o21ai_2 _06528_ (.A1(_01230_),
    .A2(_01435_),
    .B1(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__buf_1 _06529_ (.A(_01187_),
    .X(_01450_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06530_ (.A(_01244_),
    .X(_01451_));
 sky130_fd_sc_hd__nor2_2 _06531_ (.A(_01451_),
    .B(_01351_),
    .Y(_01452_));
 sky130_fd_sc_hd__a31o_2 _06532_ (.A1(_01431_),
    .A2(_01449_),
    .A3(_01450_),
    .B1(_01452_),
    .X(_01453_));
 sky130_fd_sc_hd__buf_1 _06533_ (.A(_01197_),
    .X(_01454_));
 sky130_fd_sc_hd__buf_1 _06534_ (.A(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__buf_1 _06535_ (.A(_01455_),
    .X(_01456_));
 sky130_fd_sc_hd__mux4_2 _06536_ (.A0(\rvsingle.dp.rf.rf[4][21] ),
    .A1(\rvsingle.dp.rf.rf[5][21] ),
    .A2(\rvsingle.dp.rf.rf[6][21] ),
    .A3(\rvsingle.dp.rf.rf[7][21] ),
    .S0(_01329_),
    .S1(_01456_),
    .X(_01457_));
 sky130_fd_sc_hd__nor2_2 _06537_ (.A(_01193_),
    .B(\rvsingle.dp.rf.rf[0][21] ),
    .Y(_01458_));
 sky130_fd_sc_hd__o21ai_2 _06538_ (.A1(\rvsingle.dp.rf.rf[1][21] ),
    .A2(_01441_),
    .B1(_01437_),
    .Y(_01459_));
 sky130_fd_sc_hd__buf_1 _06539_ (.A(_01206_),
    .X(_01460_));
 sky130_fd_sc_hd__buf_1 _06540_ (.A(_01460_),
    .X(_01461_));
 sky130_fd_sc_hd__buf_1 _06541_ (.A(_01190_),
    .X(_01462_));
 sky130_fd_sc_hd__buf_1 _06542_ (.A(_01462_),
    .X(_01463_));
 sky130_fd_sc_hd__o21a_2 _06543_ (.A1(_01463_),
    .A2(\rvsingle.dp.rf.rf[2][21] ),
    .B1(_01199_),
    .X(_01464_));
 sky130_fd_sc_hd__o21ai_2 _06544_ (.A1(\rvsingle.dp.rf.rf[3][21] ),
    .A2(_01296_),
    .B1(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__o211ai_2 _06545_ (.A1(_01458_),
    .A2(_01459_),
    .B1(_01461_),
    .C1(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__o211ai_2 _06546_ (.A1(_01208_),
    .A2(_01457_),
    .B1(_01466_),
    .C1(_01218_),
    .Y(_01467_));
 sky130_fd_sc_hd__buf_1 _06547_ (.A(_01190_),
    .X(_01468_));
 sky130_fd_sc_hd__buf_1 _06548_ (.A(_01468_),
    .X(_01469_));
 sky130_fd_sc_hd__buf_1 _06549_ (.A(_01454_),
    .X(_01470_));
 sky130_fd_sc_hd__buf_1 _06550_ (.A(_01470_),
    .X(_01471_));
 sky130_fd_sc_hd__mux4_2 _06551_ (.A0(\rvsingle.dp.rf.rf[8][21] ),
    .A1(\rvsingle.dp.rf.rf[9][21] ),
    .A2(\rvsingle.dp.rf.rf[10][21] ),
    .A3(\rvsingle.dp.rf.rf[11][21] ),
    .S0(_01469_),
    .S1(_01471_),
    .X(_01472_));
 sky130_fd_sc_hd__or2_2 _06552_ (.A(_01192_),
    .B(\rvsingle.dp.rf.rf[14][21] ),
    .X(_01473_));
 sky130_fd_sc_hd__o211a_2 _06553_ (.A1(_01441_),
    .A2(\rvsingle.dp.rf.rf[15][21] ),
    .B1(_01434_),
    .C1(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__or2_2 _06554_ (.A(_01192_),
    .B(\rvsingle.dp.rf.rf[12][21] ),
    .X(_01475_));
 sky130_fd_sc_hd__o211ai_2 _06555_ (.A1(\rvsingle.dp.rf.rf[13][21] ),
    .A2(_01441_),
    .B1(_01437_),
    .C1(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__nand2_2 _06556_ (.A(_01476_),
    .B(_01445_),
    .Y(_01477_));
 sky130_fd_sc_hd__buf_1 _06557_ (.A(_01446_),
    .X(_01478_));
 sky130_fd_sc_hd__o221ai_2 _06558_ (.A1(_01230_),
    .A2(_01472_),
    .B1(_01474_),
    .B2(_01477_),
    .C1(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__and3_2 _06559_ (.A(_01316_),
    .B(_01467_),
    .C(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__buf_1 _06560_ (.A(_01082_),
    .X(_01481_));
 sky130_fd_sc_hd__buf_1 _06561_ (.A(_01481_),
    .X(_01482_));
 sky130_fd_sc_hd__inv_2 _06562_ (.A(Instr[31]),
    .Y(_01483_));
 sky130_fd_sc_hd__or2_2 _06563_ (.A(_01064_),
    .B(_01073_),
    .X(_01484_));
 sky130_fd_sc_hd__buf_1 _06564_ (.A(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__buf_1 _06565_ (.A(_01485_),
    .X(_01486_));
 sky130_fd_sc_hd__buf_1 _06566_ (.A(_01086_),
    .X(_01487_));
 sky130_fd_sc_hd__buf_1 _06567_ (.A(_01487_),
    .X(_01488_));
 sky130_fd_sc_hd__buf_1 _06568_ (.A(_01103_),
    .X(_01489_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06569_ (.A(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__buf_1 _06570_ (.A(_01490_),
    .X(_01491_));
 sky130_fd_sc_hd__buf_1 _06571_ (.A(_01135_),
    .X(_01492_));
 sky130_fd_sc_hd__buf_1 _06572_ (.A(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__or2_2 _06573_ (.A(_01493_),
    .B(\rvsingle.dp.rf.rf[26][21] ),
    .X(_01494_));
 sky130_fd_sc_hd__o211a_2 _06574_ (.A1(_01488_),
    .A2(\rvsingle.dp.rf.rf[27][21] ),
    .B1(_01491_),
    .C1(_01494_),
    .X(_01495_));
 sky130_fd_sc_hd__buf_1 _06575_ (.A(_01091_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_1 _06576_ (.A(_01496_),
    .X(_01497_));
 sky130_fd_sc_hd__buf_1 _06577_ (.A(Instr[20]),
    .X(_01498_));
 sky130_fd_sc_hd__buf_1 _06578_ (.A(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__or2_2 _06579_ (.A(_01499_),
    .B(\rvsingle.dp.rf.rf[24][21] ),
    .X(_01500_));
 sky130_fd_sc_hd__or2b_2 _06580_ (.A(\rvsingle.dp.rf.rf[25][21] ),
    .B_N(_01493_),
    .X(_01501_));
 sky130_fd_sc_hd__buf_1 _06581_ (.A(_01110_),
    .X(_01502_));
 sky130_fd_sc_hd__buf_1 _06582_ (.A(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__a31o_2 _06583_ (.A1(_01497_),
    .A2(_01500_),
    .A3(_01501_),
    .B1(_01503_),
    .X(_01504_));
 sky130_fd_sc_hd__buf_1 _06584_ (.A(_01115_),
    .X(_01505_));
 sky130_fd_sc_hd__buf_1 _06585_ (.A(_01505_),
    .X(_01506_));
 sky130_fd_sc_hd__nor2_2 _06586_ (.A(_01269_),
    .B(\rvsingle.dp.rf.rf[30][21] ),
    .Y(_01507_));
 sky130_fd_sc_hd__buf_1 _06587_ (.A(_01086_),
    .X(_01508_));
 sky130_fd_sc_hd__buf_1 _06588_ (.A(_01508_),
    .X(_01509_));
 sky130_fd_sc_hd__o21ai_2 _06589_ (.A1(\rvsingle.dp.rf.rf[31][21] ),
    .A2(_01509_),
    .B1(_01491_),
    .Y(_01510_));
 sky130_fd_sc_hd__buf_1 _06590_ (.A(_01110_),
    .X(_01511_));
 sky130_fd_sc_hd__buf_1 _06591_ (.A(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__buf_1 _06592_ (.A(_01267_),
    .X(_01513_));
 sky130_fd_sc_hd__or2_2 _06593_ (.A(_01513_),
    .B(\rvsingle.dp.rf.rf[28][21] ),
    .X(_01514_));
 sky130_fd_sc_hd__o211ai_2 _06594_ (.A1(\rvsingle.dp.rf.rf[29][21] ),
    .A2(_01488_),
    .B1(_01497_),
    .C1(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__o211ai_2 _06595_ (.A1(_01507_),
    .A2(_01510_),
    .B1(_01512_),
    .C1(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__o211ai_2 _06596_ (.A1(_01495_),
    .A2(_01504_),
    .B1(_01506_),
    .C1(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__buf_1 _06597_ (.A(_01136_),
    .X(_01518_));
 sky130_fd_sc_hd__buf_1 _06598_ (.A(_01103_),
    .X(_01519_));
 sky130_fd_sc_hd__buf_1 _06599_ (.A(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__o21ba_2 _06600_ (.A1(_01518_),
    .A2(\rvsingle.dp.rf.rf[20][21] ),
    .B1_N(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__o21ai_2 _06601_ (.A1(_01509_),
    .A2(\rvsingle.dp.rf.rf[21][21] ),
    .B1(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__buf_1 _06602_ (.A(_01489_),
    .X(_01523_));
 sky130_fd_sc_hd__o21a_2 _06603_ (.A1(_01493_),
    .A2(\rvsingle.dp.rf.rf[22][21] ),
    .B1(_01523_),
    .X(_01524_));
 sky130_fd_sc_hd__o21ai_2 _06604_ (.A1(\rvsingle.dp.rf.rf[23][21] ),
    .A2(_01509_),
    .B1(_01524_),
    .Y(_01525_));
 sky130_fd_sc_hd__buf_1 _06605_ (.A(_01115_),
    .X(_01526_));
 sky130_fd_sc_hd__a31oi_2 _06606_ (.A1(_01522_),
    .A2(_01112_),
    .A3(_01525_),
    .B1(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_2 _06607_ (.A(_01269_),
    .B(\rvsingle.dp.rf.rf[16][21] ),
    .Y(_01528_));
 sky130_fd_sc_hd__o21ai_2 _06608_ (.A1(\rvsingle.dp.rf.rf[17][21] ),
    .A2(_01509_),
    .B1(_01497_),
    .Y(_01529_));
 sky130_fd_sc_hd__dlymetal6s4s_1 _06609_ (.A(_01103_),
    .X(_01530_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _06610_ (.A(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__o21a_2 _06611_ (.A1(_01256_),
    .A2(\rvsingle.dp.rf.rf[18][21] ),
    .B1(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__o21ai_2 _06612_ (.A1(\rvsingle.dp.rf.rf[19][21] ),
    .A2(_01488_),
    .B1(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__o211ai_2 _06613_ (.A1(_01528_),
    .A2(_01529_),
    .B1(_01132_),
    .C1(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__nand2_2 _06614_ (.A(_01527_),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__nand3_2 _06615_ (.A(_01517_),
    .B(_01535_),
    .C(_01147_),
    .Y(_01536_));
 sky130_fd_sc_hd__buf_1 _06616_ (.A(_01083_),
    .X(_01537_));
 sky130_fd_sc_hd__nor2_2 _06617_ (.A(_01383_),
    .B(\rvsingle.dp.rf.rf[14][21] ),
    .Y(_01538_));
 sky130_fd_sc_hd__buf_1 _06618_ (.A(_01086_),
    .X(_01539_));
 sky130_fd_sc_hd__buf_1 _06619_ (.A(_01539_),
    .X(_01540_));
 sky130_fd_sc_hd__o21ai_2 _06620_ (.A1(\rvsingle.dp.rf.rf[15][21] ),
    .A2(_01540_),
    .B1(_01260_),
    .Y(_01541_));
 sky130_fd_sc_hd__buf_1 _06621_ (.A(_01091_),
    .X(_01542_));
 sky130_fd_sc_hd__buf_1 _06622_ (.A(_01542_),
    .X(_01543_));
 sky130_fd_sc_hd__buf_1 _06623_ (.A(_01095_),
    .X(_01544_));
 sky130_fd_sc_hd__buf_1 _06624_ (.A(_01544_),
    .X(_01545_));
 sky130_fd_sc_hd__or2_2 _06625_ (.A(_01545_),
    .B(\rvsingle.dp.rf.rf[12][21] ),
    .X(_01546_));
 sky130_fd_sc_hd__o211ai_2 _06626_ (.A1(\rvsingle.dp.rf.rf[13][21] ),
    .A2(_01540_),
    .B1(_01543_),
    .C1(_01546_),
    .Y(_01547_));
 sky130_fd_sc_hd__o211ai_2 _06627_ (.A1(_01538_),
    .A2(_01541_),
    .B1(_01547_),
    .C1(_01512_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_2 _06628_ (.A(_01383_),
    .B(\rvsingle.dp.rf.rf[8][21] ),
    .Y(_01549_));
 sky130_fd_sc_hd__o21ai_2 _06629_ (.A1(\rvsingle.dp.rf.rf[9][21] ),
    .A2(_01540_),
    .B1(_01543_),
    .Y(_01550_));
 sky130_fd_sc_hd__buf_1 _06630_ (.A(_01103_),
    .X(_01551_));
 sky130_fd_sc_hd__buf_1 _06631_ (.A(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__o21a_2 _06632_ (.A1(_01137_),
    .A2(\rvsingle.dp.rf.rf[10][21] ),
    .B1(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__o21ai_2 _06633_ (.A1(\rvsingle.dp.rf.rf[11][21] ),
    .A2(_01509_),
    .B1(_01553_),
    .Y(_01554_));
 sky130_fd_sc_hd__o211ai_2 _06634_ (.A1(_01549_),
    .A2(_01550_),
    .B1(_01132_),
    .C1(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand3_2 _06635_ (.A(_01548_),
    .B(_01555_),
    .C(_01506_),
    .Y(_01556_));
 sky130_fd_sc_hd__buf_1 _06636_ (.A(_01095_),
    .X(_01557_));
 sky130_fd_sc_hd__buf_1 _06637_ (.A(_01557_),
    .X(_01558_));
 sky130_fd_sc_hd__buf_1 _06638_ (.A(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__nor2_2 _06639_ (.A(_01559_),
    .B(\rvsingle.dp.rf.rf[0][21] ),
    .Y(_01560_));
 sky130_fd_sc_hd__buf_1 _06640_ (.A(_01135_),
    .X(_01561_));
 sky130_fd_sc_hd__buf_1 _06641_ (.A(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__and2b_2 _06642_ (.A_N(\rvsingle.dp.rf.rf[1][21] ),
    .B(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__buf_1 _06643_ (.A(_01130_),
    .X(_01564_));
 sky130_fd_sc_hd__buf_1 _06644_ (.A(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__buf_1 _06645_ (.A(_01095_),
    .X(_01566_));
 sky130_fd_sc_hd__buf_1 _06646_ (.A(_01566_),
    .X(_01567_));
 sky130_fd_sc_hd__or2b_2 _06647_ (.A(\rvsingle.dp.rf.rf[3][21] ),
    .B_N(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__o211ai_2 _06648_ (.A1(_01559_),
    .A2(\rvsingle.dp.rf.rf[2][21] ),
    .B1(_01260_),
    .C1(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__o311ai_2 _06649_ (.A1(_01491_),
    .A2(_01560_),
    .A3(_01563_),
    .B1(_01565_),
    .C1(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__nor2_2 _06650_ (.A(_01559_),
    .B(\rvsingle.dp.rf.rf[6][21] ),
    .Y(_01571_));
 sky130_fd_sc_hd__and2b_2 _06651_ (.A_N(\rvsingle.dp.rf.rf[7][21] ),
    .B(_01562_),
    .X(_01572_));
 sky130_fd_sc_hd__o21ba_2 _06652_ (.A1(_01499_),
    .A2(\rvsingle.dp.rf.rf[4][21] ),
    .B1_N(_01259_),
    .X(_01573_));
 sky130_fd_sc_hd__o21ai_2 _06653_ (.A1(_01540_),
    .A2(\rvsingle.dp.rf.rf[5][21] ),
    .B1(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__o311ai_2 _06654_ (.A1(_01497_),
    .A2(_01571_),
    .A3(_01572_),
    .B1(_01112_),
    .C1(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__nand3_2 _06655_ (.A(_01157_),
    .B(_01570_),
    .C(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__nand3_2 _06656_ (.A(_01378_),
    .B(_01556_),
    .C(_01576_),
    .Y(_01577_));
 sky130_fd_sc_hd__nand4_2 _06657_ (.A(_01536_),
    .B(_01537_),
    .C(_01153_),
    .D(_01577_),
    .Y(_01578_));
 sky130_fd_sc_hd__o211a_2 _06658_ (.A1(_01482_),
    .A2(_01483_),
    .B1(_01486_),
    .C1(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__o21ai_2 _06659_ (.A1(_01171_),
    .A2(_01176_),
    .B1(_01177_),
    .Y(_01580_));
 sky130_fd_sc_hd__buf_1 _06660_ (.A(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__a21oi_2 _06661_ (.A1(_01581_),
    .A2(_01578_),
    .B1(_01486_),
    .Y(_01582_));
 sky130_fd_sc_hd__o22ai_2 _06662_ (.A1(_01453_),
    .A2(_01480_),
    .B1(_01579_),
    .B2(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__buf_1 _06663_ (.A(_01183_),
    .X(_01584_));
 sky130_fd_sc_hd__a41o_2 _06664_ (.A1(_01153_),
    .A2(_01536_),
    .A3(_01577_),
    .A4(_01482_),
    .B1(_01584_),
    .X(_01585_));
 sky130_fd_sc_hd__nor2_2 _06665_ (.A(_01480_),
    .B(_01453_),
    .Y(_01586_));
 sky130_fd_sc_hd__buf_1 _06666_ (.A(_01580_),
    .X(_01587_));
 sky130_fd_sc_hd__a21o_2 _06667_ (.A1(_01587_),
    .A2(_01578_),
    .B1(_01486_),
    .X(_01588_));
 sky130_fd_sc_hd__o211ai_2 _06668_ (.A1(_01179_),
    .A2(_01585_),
    .B1(_01586_),
    .C1(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__nand2_2 _06669_ (.A(_01583_),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__buf_1 _06670_ (.A(_01485_),
    .X(_01591_));
 sky130_fd_sc_hd__buf_1 _06671_ (.A(_01152_),
    .X(_01592_));
 sky130_fd_sc_hd__buf_1 _06672_ (.A(_01376_),
    .X(_01593_));
 sky130_fd_sc_hd__buf_1 _06673_ (.A(_01095_),
    .X(_01594_));
 sky130_fd_sc_hd__buf_1 _06674_ (.A(_01594_),
    .X(_01595_));
 sky130_fd_sc_hd__buf_1 _06675_ (.A(_01103_),
    .X(_01596_));
 sky130_fd_sc_hd__o21bai_2 _06676_ (.A1(_01595_),
    .A2(\rvsingle.dp.rf.rf[8][20] ),
    .B1_N(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__and2b_2 _06677_ (.A_N(\rvsingle.dp.rf.rf[9][20] ),
    .B(_01097_),
    .X(_01598_));
 sky130_fd_sc_hd__buf_1 _06678_ (.A(_01130_),
    .X(_01599_));
 sky130_fd_sc_hd__buf_1 _06679_ (.A(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__o21ai_2 _06680_ (.A1(_01597_),
    .A2(_01598_),
    .B1(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__buf_1 _06681_ (.A(_01135_),
    .X(_01602_));
 sky130_fd_sc_hd__buf_1 _06682_ (.A(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__buf_1 _06683_ (.A(_01103_),
    .X(_01604_));
 sky130_fd_sc_hd__buf_1 _06684_ (.A(_01604_),
    .X(_01605_));
 sky130_fd_sc_hd__buf_1 _06685_ (.A(Instr[20]),
    .X(_01606_));
 sky130_fd_sc_hd__buf_1 _06686_ (.A(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__or2b_2 _06687_ (.A(\rvsingle.dp.rf.rf[11][20] ),
    .B_N(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__o211a_2 _06688_ (.A1(_01603_),
    .A2(\rvsingle.dp.rf.rf[10][20] ),
    .B1(_01605_),
    .C1(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__buf_1 _06689_ (.A(Instr[21]),
    .X(_01610_));
 sky130_fd_sc_hd__buf_1 _06690_ (.A(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__buf_1 _06691_ (.A(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__buf_1 _06692_ (.A(_01095_),
    .X(_01613_));
 sky130_fd_sc_hd__buf_1 _06693_ (.A(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__nor2_2 _06694_ (.A(_01614_),
    .B(\rvsingle.dp.rf.rf[12][20] ),
    .Y(_01615_));
 sky130_fd_sc_hd__and2b_2 _06695_ (.A_N(\rvsingle.dp.rf.rf[13][20] ),
    .B(_01148_),
    .X(_01616_));
 sky130_fd_sc_hd__buf_1 _06696_ (.A(_01110_),
    .X(_01617_));
 sky130_fd_sc_hd__buf_1 _06697_ (.A(_01135_),
    .X(_01618_));
 sky130_fd_sc_hd__buf_1 _06698_ (.A(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__buf_1 _06699_ (.A(_01530_),
    .X(_01620_));
 sky130_fd_sc_hd__or2b_2 _06700_ (.A(\rvsingle.dp.rf.rf[15][20] ),
    .B_N(_01255_),
    .X(_01621_));
 sky130_fd_sc_hd__o211ai_2 _06701_ (.A1(_01619_),
    .A2(\rvsingle.dp.rf.rf[14][20] ),
    .B1(_01620_),
    .C1(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__o311ai_2 _06702_ (.A1(_01612_),
    .A2(_01615_),
    .A3(_01616_),
    .B1(_01617_),
    .C1(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__o211ai_2 _06703_ (.A1(_01601_),
    .A2(_01609_),
    .B1(_01116_),
    .C1(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__inv_2 _06704_ (.A(\rvsingle.dp.rf.rf[5][20] ),
    .Y(_01625_));
 sky130_fd_sc_hd__buf_1 _06705_ (.A(_01611_),
    .X(_01626_));
 sky130_fd_sc_hd__nor2_2 _06706_ (.A(_01256_),
    .B(\rvsingle.dp.rf.rf[4][20] ),
    .Y(_01627_));
 sky130_fd_sc_hd__a211oi_2 _06707_ (.A1(_01625_),
    .A2(_01098_),
    .B1(_01626_),
    .C1(_01627_),
    .Y(_01628_));
 sky130_fd_sc_hd__o21ai_2 _06708_ (.A1(_01518_),
    .A2(\rvsingle.dp.rf.rf[6][20] ),
    .B1(_01620_),
    .Y(_01629_));
 sky130_fd_sc_hd__buf_1 _06709_ (.A(_01557_),
    .X(_01630_));
 sky130_fd_sc_hd__and2b_2 _06710_ (.A_N(\rvsingle.dp.rf.rf[7][20] ),
    .B(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__buf_1 _06711_ (.A(_01110_),
    .X(_01632_));
 sky130_fd_sc_hd__o21ai_2 _06712_ (.A1(_01629_),
    .A2(_01631_),
    .B1(_01632_),
    .Y(_01633_));
 sky130_fd_sc_hd__buf_1 _06713_ (.A(_01155_),
    .X(_01634_));
 sky130_fd_sc_hd__nor2_2 _06714_ (.A(_01614_),
    .B(\rvsingle.dp.rf.rf[0][20] ),
    .Y(_01635_));
 sky130_fd_sc_hd__and2b_2 _06715_ (.A_N(\rvsingle.dp.rf.rf[1][20] ),
    .B(_01148_),
    .X(_01636_));
 sky130_fd_sc_hd__or2b_2 _06716_ (.A(\rvsingle.dp.rf.rf[3][20] ),
    .B_N(_01255_),
    .X(_01637_));
 sky130_fd_sc_hd__o211ai_2 _06717_ (.A1(_01619_),
    .A2(\rvsingle.dp.rf.rf[2][20] ),
    .B1(_01620_),
    .C1(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__o311ai_2 _06718_ (.A1(_01612_),
    .A2(_01635_),
    .A3(_01636_),
    .B1(_01600_),
    .C1(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__o211ai_2 _06719_ (.A1(_01628_),
    .A2(_01633_),
    .B1(_01634_),
    .C1(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__nand3_2 _06720_ (.A(_01593_),
    .B(_01624_),
    .C(_01640_),
    .Y(_01641_));
 sky130_fd_sc_hd__buf_1 _06721_ (.A(_01606_),
    .X(_01642_));
 sky130_fd_sc_hd__buf_1 _06722_ (.A(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__nor2_2 _06723_ (.A(_01643_),
    .B(\rvsingle.dp.rf.rf[30][20] ),
    .Y(_01644_));
 sky130_fd_sc_hd__buf_1 _06724_ (.A(_01086_),
    .X(_01645_));
 sky130_fd_sc_hd__buf_1 _06725_ (.A(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__buf_1 _06726_ (.A(_01103_),
    .X(_01647_));
 sky130_fd_sc_hd__buf_1 _06727_ (.A(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__o21ai_2 _06728_ (.A1(\rvsingle.dp.rf.rf[31][20] ),
    .A2(_01646_),
    .B1(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__buf_1 _06729_ (.A(_01135_),
    .X(_01650_));
 sky130_fd_sc_hd__or2_2 _06730_ (.A(_01650_),
    .B(\rvsingle.dp.rf.rf[28][20] ),
    .X(_01651_));
 sky130_fd_sc_hd__o211ai_2 _06731_ (.A1(\rvsingle.dp.rf.rf[29][20] ),
    .A2(_01646_),
    .B1(_01092_),
    .C1(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__o211ai_2 _06732_ (.A1(_01644_),
    .A2(_01649_),
    .B1(_01652_),
    .C1(_01503_),
    .Y(_01653_));
 sky130_fd_sc_hd__buf_1 _06733_ (.A(_01610_),
    .X(_01654_));
 sky130_fd_sc_hd__buf_1 _06734_ (.A(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__buf_1 _06735_ (.A(_01561_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_2 _06736_ (.A(_01656_),
    .B(\rvsingle.dp.rf.rf[24][20] ),
    .Y(_01657_));
 sky130_fd_sc_hd__buf_1 _06737_ (.A(_01557_),
    .X(_01658_));
 sky130_fd_sc_hd__and2b_2 _06738_ (.A_N(\rvsingle.dp.rf.rf[25][20] ),
    .B(_01658_),
    .X(_01659_));
 sky130_fd_sc_hd__buf_1 _06739_ (.A(_01604_),
    .X(_01660_));
 sky130_fd_sc_hd__or2b_2 _06740_ (.A(\rvsingle.dp.rf.rf[27][20] ),
    .B_N(_01602_),
    .X(_01661_));
 sky130_fd_sc_hd__o211ai_2 _06741_ (.A1(_01656_),
    .A2(\rvsingle.dp.rf.rf[26][20] ),
    .B1(_01660_),
    .C1(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__o311ai_2 _06742_ (.A1(_01655_),
    .A2(_01657_),
    .A3(_01659_),
    .B1(_01600_),
    .C1(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__nand3_2 _06743_ (.A(_01653_),
    .B(_01663_),
    .C(_01526_),
    .Y(_01664_));
 sky130_fd_sc_hd__inv_2 _06744_ (.A(\rvsingle.dp.rf.rf[23][20] ),
    .Y(_01665_));
 sky130_fd_sc_hd__buf_1 _06745_ (.A(_01148_),
    .X(_01666_));
 sky130_fd_sc_hd__buf_1 _06746_ (.A(_01091_),
    .X(_01667_));
 sky130_fd_sc_hd__buf_1 _06747_ (.A(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__nor2_2 _06748_ (.A(_01256_),
    .B(\rvsingle.dp.rf.rf[22][20] ),
    .Y(_01669_));
 sky130_fd_sc_hd__a211oi_2 _06749_ (.A1(_01665_),
    .A2(_01666_),
    .B1(_01668_),
    .C1(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__o21bai_2 _06750_ (.A1(_01137_),
    .A2(\rvsingle.dp.rf.rf[20][20] ),
    .B1_N(_01611_),
    .Y(_01671_));
 sky130_fd_sc_hd__and2b_2 _06751_ (.A_N(\rvsingle.dp.rf.rf[21][20] ),
    .B(_01558_),
    .X(_01672_));
 sky130_fd_sc_hd__o21ai_2 _06752_ (.A1(_01671_),
    .A2(_01672_),
    .B1(_01617_),
    .Y(_01673_));
 sky130_fd_sc_hd__nor2_2 _06753_ (.A(_01614_),
    .B(\rvsingle.dp.rf.rf[18][20] ),
    .Y(_01674_));
 sky130_fd_sc_hd__buf_1 _06754_ (.A(_01096_),
    .X(_01675_));
 sky130_fd_sc_hd__and2b_2 _06755_ (.A_N(\rvsingle.dp.rf.rf[19][20] ),
    .B(_01675_),
    .X(_01676_));
 sky130_fd_sc_hd__buf_1 _06756_ (.A(_01645_),
    .X(_01677_));
 sky130_fd_sc_hd__o21ba_2 _06757_ (.A1(_01602_),
    .A2(\rvsingle.dp.rf.rf[16][20] ),
    .B1_N(_01551_),
    .X(_01678_));
 sky130_fd_sc_hd__o21ai_2 _06758_ (.A1(_01677_),
    .A2(\rvsingle.dp.rf.rf[17][20] ),
    .B1(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__o311ai_2 _06759_ (.A1(_01092_),
    .A2(_01674_),
    .A3(_01676_),
    .B1(_01679_),
    .C1(_01600_),
    .Y(_01680_));
 sky130_fd_sc_hd__o211ai_2 _06760_ (.A1(_01670_),
    .A2(_01673_),
    .B1(_01634_),
    .C1(_01680_),
    .Y(_01681_));
 sky130_fd_sc_hd__buf_1 _06761_ (.A(_01145_),
    .X(_01682_));
 sky130_fd_sc_hd__nand3_2 _06762_ (.A(_01664_),
    .B(_01681_),
    .C(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand4_2 _06763_ (.A(_01592_),
    .B(_01641_),
    .C(_01683_),
    .D(_01481_),
    .Y(_01684_));
 sky130_fd_sc_hd__o211a_2 _06764_ (.A1(_01084_),
    .A2(_01483_),
    .B1(_01591_),
    .C1(_01684_),
    .X(_01685_));
 sky130_fd_sc_hd__mux4_2 _06765_ (.A0(\rvsingle.dp.rf.rf[8][20] ),
    .A1(\rvsingle.dp.rf.rf[9][20] ),
    .A2(\rvsingle.dp.rf.rf[10][20] ),
    .A3(\rvsingle.dp.rf.rf[11][20] ),
    .S0(_01463_),
    .S1(_01471_),
    .X(_01686_));
 sky130_fd_sc_hd__buf_1 _06766_ (.A(_01293_),
    .X(_01687_));
 sky130_fd_sc_hd__buf_1 _06767_ (.A(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__buf_1 _06768_ (.A(_01307_),
    .X(_01689_));
 sky130_fd_sc_hd__buf_1 _06769_ (.A(_01190_),
    .X(_01690_));
 sky130_fd_sc_hd__buf_1 _06770_ (.A(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__or2_2 _06771_ (.A(_01691_),
    .B(\rvsingle.dp.rf.rf[12][20] ),
    .X(_01692_));
 sky130_fd_sc_hd__o211ai_2 _06772_ (.A1(\rvsingle.dp.rf.rf[13][20] ),
    .A2(_01688_),
    .B1(_01689_),
    .C1(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__buf_1 _06773_ (.A(_01444_),
    .X(_01694_));
 sky130_fd_sc_hd__buf_1 _06774_ (.A(_01349_),
    .X(_01695_));
 sky130_fd_sc_hd__buf_1 _06775_ (.A(_01299_),
    .X(_01696_));
 sky130_fd_sc_hd__o21a_2 _06776_ (.A1(_01695_),
    .A2(\rvsingle.dp.rf.rf[14][20] ),
    .B1(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__o21ai_2 _06777_ (.A1(\rvsingle.dp.rf.rf[15][20] ),
    .A2(_01688_),
    .B1(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__buf_1 _06778_ (.A(_01216_),
    .X(_01699_));
 sky130_fd_sc_hd__a31oi_2 _06779_ (.A1(_01693_),
    .A2(_01694_),
    .A3(_01698_),
    .B1(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__o21ai_2 _06780_ (.A1(_01230_),
    .A2(_01686_),
    .B1(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__buf_1 _06781_ (.A(_01172_),
    .X(_01702_));
 sky130_fd_sc_hd__buf_1 _06782_ (.A(_01702_),
    .X(_01703_));
 sky130_fd_sc_hd__mux4_2 _06783_ (.A0(\rvsingle.dp.rf.rf[0][20] ),
    .A1(\rvsingle.dp.rf.rf[1][20] ),
    .A2(\rvsingle.dp.rf.rf[2][20] ),
    .A3(\rvsingle.dp.rf.rf[3][20] ),
    .S0(_01469_),
    .S1(_01471_),
    .X(_01704_));
 sky130_fd_sc_hd__nor2_2 _06784_ (.A(_01420_),
    .B(\rvsingle.dp.rf.rf[4][20] ),
    .Y(_01705_));
 sky130_fd_sc_hd__a211o_2 _06785_ (.A1(_01625_),
    .A2(_01329_),
    .B1(_01199_),
    .C1(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__buf_1 _06786_ (.A(_01419_),
    .X(_01707_));
 sky130_fd_sc_hd__buf_1 _06787_ (.A(_01454_),
    .X(_01708_));
 sky130_fd_sc_hd__o21a_2 _06788_ (.A1(_01707_),
    .A2(\rvsingle.dp.rf.rf[6][20] ),
    .B1(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__o21ai_2 _06789_ (.A1(\rvsingle.dp.rf.rf[7][20] ),
    .A2(_01688_),
    .B1(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__buf_1 _06790_ (.A(_01444_),
    .X(_01711_));
 sky130_fd_sc_hd__a31oi_2 _06791_ (.A1(_01706_),
    .A2(_01710_),
    .A3(_01711_),
    .B1(_01221_),
    .Y(_01712_));
 sky130_fd_sc_hd__o21ai_2 _06792_ (.A1(_01703_),
    .A2(_01704_),
    .B1(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__nand2_2 _06793_ (.A(_01701_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__mux2_2 _06794_ (.A0(\rvsingle.dp.rf.rf[16][20] ),
    .A1(\rvsingle.dp.rf.rf[17][20] ),
    .S(_01417_),
    .X(_01715_));
 sky130_fd_sc_hd__buf_1 _06795_ (.A(_01307_),
    .X(_01716_));
 sky130_fd_sc_hd__buf_1 _06796_ (.A(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__or2_2 _06797_ (.A(_01707_),
    .B(\rvsingle.dp.rf.rf[18][20] ),
    .X(_01718_));
 sky130_fd_sc_hd__o211a_2 _06798_ (.A1(_01688_),
    .A2(\rvsingle.dp.rf.rf[19][20] ),
    .B1(_01456_),
    .C1(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__a211oi_2 _06799_ (.A1(_01715_),
    .A2(_01717_),
    .B1(_01703_),
    .C1(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__buf_1 _06800_ (.A(_01206_),
    .X(_01721_));
 sky130_fd_sc_hd__buf_1 _06801_ (.A(_01721_),
    .X(_01722_));
 sky130_fd_sc_hd__mux4_2 _06802_ (.A0(\rvsingle.dp.rf.rf[20][20] ),
    .A1(\rvsingle.dp.rf.rf[21][20] ),
    .A2(\rvsingle.dp.rf.rf[22][20] ),
    .A3(\rvsingle.dp.rf.rf[23][20] ),
    .S0(_01192_),
    .S1(_01244_),
    .X(_01723_));
 sky130_fd_sc_hd__o21ai_2 _06803_ (.A1(_01722_),
    .A2(_01723_),
    .B1(_01218_),
    .Y(_01724_));
 sky130_fd_sc_hd__buf_1 _06804_ (.A(_01190_),
    .X(_01725_));
 sky130_fd_sc_hd__buf_1 _06805_ (.A(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__buf_1 _06806_ (.A(_01197_),
    .X(_01727_));
 sky130_fd_sc_hd__buf_1 _06807_ (.A(_01727_),
    .X(_01728_));
 sky130_fd_sc_hd__mux4_2 _06808_ (.A0(\rvsingle.dp.rf.rf[24][20] ),
    .A1(\rvsingle.dp.rf.rf[25][20] ),
    .A2(\rvsingle.dp.rf.rf[26][20] ),
    .A3(\rvsingle.dp.rf.rf[27][20] ),
    .S0(_01726_),
    .S1(_01728_),
    .X(_01729_));
 sky130_fd_sc_hd__buf_1 _06809_ (.A(_01425_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_2 _06810_ (.A0(\rvsingle.dp.rf.rf[28][20] ),
    .A1(\rvsingle.dp.rf.rf[29][20] ),
    .S(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__o21a_2 _06811_ (.A1(_01462_),
    .A2(\rvsingle.dp.rf.rf[30][20] ),
    .B1(_01198_),
    .X(_01732_));
 sky130_fd_sc_hd__o21a_2 _06812_ (.A1(_01295_),
    .A2(\rvsingle.dp.rf.rf[31][20] ),
    .B1(_01732_),
    .X(_01733_));
 sky130_fd_sc_hd__a211o_2 _06813_ (.A1(_01731_),
    .A2(_01437_),
    .B1(_01721_),
    .C1(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__o211ai_2 _06814_ (.A1(_01703_),
    .A2(_01729_),
    .B1(_01734_),
    .C1(_01478_),
    .Y(_01735_));
 sky130_fd_sc_hd__o211ai_2 _06815_ (.A1(_01720_),
    .A2(_01724_),
    .B1(_01188_),
    .C1(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__o211a_2 _06816_ (.A1(_01450_),
    .A2(_01714_),
    .B1(_01736_),
    .C1(_01247_),
    .X(_01737_));
 sky130_fd_sc_hd__a21o_2 _06817_ (.A1(_01587_),
    .A2(_01684_),
    .B1(_01486_),
    .X(_01738_));
 sky130_fd_sc_hd__nand3b_2 _06818_ (.A_N(_01685_),
    .B(_01737_),
    .C(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__a21oi_2 _06819_ (.A1(_01581_),
    .A2(_01684_),
    .B1(_01486_),
    .Y(_01740_));
 sky130_fd_sc_hd__o21bai_2 _06820_ (.A1(_01740_),
    .A2(_01685_),
    .B1_N(_01737_),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_2 _06821_ (.A(_01739_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__buf_1 _06822_ (.A(_01124_),
    .X(_01743_));
 sky130_fd_sc_hd__buf_1 _06823_ (.A(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__nor2_2 _06824_ (.A(_01744_),
    .B(\rvsingle.dp.rf.rf[12][23] ),
    .Y(_01745_));
 sky130_fd_sc_hd__o21bai_2 _06825_ (.A1(\rvsingle.dp.rf.rf[13][23] ),
    .A2(_01646_),
    .B1_N(_01520_),
    .Y(_01746_));
 sky130_fd_sc_hd__or2_2 _06826_ (.A(_01125_),
    .B(\rvsingle.dp.rf.rf[14][23] ),
    .X(_01747_));
 sky130_fd_sc_hd__o211ai_2 _06827_ (.A1(_01646_),
    .A2(\rvsingle.dp.rf.rf[15][23] ),
    .B1(_01105_),
    .C1(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__o211ai_2 _06828_ (.A1(_01745_),
    .A2(_01746_),
    .B1(_01632_),
    .C1(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__or2b_2 _06829_ (.A(\rvsingle.dp.rf.rf[11][23] ),
    .B_N(_01125_),
    .X(_01750_));
 sky130_fd_sc_hd__o211ai_2 _06830_ (.A1(_01603_),
    .A2(\rvsingle.dp.rf.rf[10][23] ),
    .B1(_01605_),
    .C1(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__buf_1 _06831_ (.A(Instr[20]),
    .X(_01752_));
 sky130_fd_sc_hd__buf_1 _06832_ (.A(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__o21ba_2 _06833_ (.A1(_01753_),
    .A2(\rvsingle.dp.rf.rf[8][23] ),
    .B1_N(_01604_),
    .X(_01754_));
 sky130_fd_sc_hd__o21ai_2 _06834_ (.A1(_01646_),
    .A2(\rvsingle.dp.rf.rf[9][23] ),
    .B1(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__nand3_2 _06835_ (.A(_01565_),
    .B(_01751_),
    .C(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__nand3_2 _06836_ (.A(_01749_),
    .B(_01756_),
    .C(_01526_),
    .Y(_01757_));
 sky130_fd_sc_hd__inv_2 _06837_ (.A(\rvsingle.dp.rf.rf[7][23] ),
    .Y(_01758_));
 sky130_fd_sc_hd__buf_1 _06838_ (.A(_01667_),
    .X(_01759_));
 sky130_fd_sc_hd__nor2_2 _06839_ (.A(_01603_),
    .B(\rvsingle.dp.rf.rf[6][23] ),
    .Y(_01760_));
 sky130_fd_sc_hd__a211oi_2 _06840_ (.A1(_01758_),
    .A2(_01559_),
    .B1(_01759_),
    .C1(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__o21bai_2 _06841_ (.A1(_01619_),
    .A2(\rvsingle.dp.rf.rf[4][23] ),
    .B1_N(_01654_),
    .Y(_01762_));
 sky130_fd_sc_hd__buf_1 _06842_ (.A(_01381_),
    .X(_01763_));
 sky130_fd_sc_hd__and2b_2 _06843_ (.A_N(\rvsingle.dp.rf.rf[5][23] ),
    .B(_01763_),
    .X(_01764_));
 sky130_fd_sc_hd__o21ai_2 _06844_ (.A1(_01762_),
    .A2(_01764_),
    .B1(_01632_),
    .Y(_01765_));
 sky130_fd_sc_hd__nor2_2 _06845_ (.A(_01656_),
    .B(\rvsingle.dp.rf.rf[0][23] ),
    .Y(_01766_));
 sky130_fd_sc_hd__and2b_2 _06846_ (.A_N(\rvsingle.dp.rf.rf[1][23] ),
    .B(_01658_),
    .X(_01767_));
 sky130_fd_sc_hd__buf_1 _06847_ (.A(_01599_),
    .X(_01768_));
 sky130_fd_sc_hd__buf_1 _06848_ (.A(_01135_),
    .X(_01769_));
 sky130_fd_sc_hd__or2b_2 _06849_ (.A(\rvsingle.dp.rf.rf[3][23] ),
    .B_N(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__o211ai_2 _06850_ (.A1(_01656_),
    .A2(\rvsingle.dp.rf.rf[2][23] ),
    .B1(_01660_),
    .C1(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__o311ai_2 _06851_ (.A1(_01655_),
    .A2(_01766_),
    .A3(_01767_),
    .B1(_01768_),
    .C1(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__o211ai_2 _06852_ (.A1(_01761_),
    .A2(_01765_),
    .B1(_01634_),
    .C1(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__nand3_2 _06853_ (.A(_01593_),
    .B(_01757_),
    .C(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hd__or2b_2 _06854_ (.A(\rvsingle.dp.rf.rf[27][23] ),
    .B_N(_01753_),
    .X(_01775_));
 sky130_fd_sc_hd__o211a_2 _06855_ (.A1(_01744_),
    .A2(\rvsingle.dp.rf.rf[26][23] ),
    .B1(_01648_),
    .C1(_01775_),
    .X(_01776_));
 sky130_fd_sc_hd__buf_1 _06856_ (.A(_01258_),
    .X(_01777_));
 sky130_fd_sc_hd__o21bai_2 _06857_ (.A1(_01656_),
    .A2(\rvsingle.dp.rf.rf[24][23] ),
    .B1_N(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__buf_1 _06858_ (.A(_01095_),
    .X(_01779_));
 sky130_fd_sc_hd__buf_1 _06859_ (.A(_01779_),
    .X(_01780_));
 sky130_fd_sc_hd__and2b_2 _06860_ (.A_N(\rvsingle.dp.rf.rf[25][23] ),
    .B(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__o21ai_2 _06861_ (.A1(_01778_),
    .A2(_01781_),
    .B1(_01768_),
    .Y(_01782_));
 sky130_fd_sc_hd__nor2_2 _06862_ (.A(_01643_),
    .B(\rvsingle.dp.rf.rf[28][23] ),
    .Y(_01783_));
 sky130_fd_sc_hd__o21bai_2 _06863_ (.A1(\rvsingle.dp.rf.rf[29][23] ),
    .A2(_01646_),
    .B1_N(_01520_),
    .Y(_01784_));
 sky130_fd_sc_hd__or2_2 _06864_ (.A(_01125_),
    .B(\rvsingle.dp.rf.rf[30][23] ),
    .X(_01785_));
 sky130_fd_sc_hd__o211ai_2 _06865_ (.A1(_01646_),
    .A2(\rvsingle.dp.rf.rf[31][23] ),
    .B1(_01648_),
    .C1(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__o211ai_2 _06866_ (.A1(_01783_),
    .A2(_01784_),
    .B1(_01632_),
    .C1(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__o211ai_2 _06867_ (.A1(_01776_),
    .A2(_01782_),
    .B1(_01526_),
    .C1(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__o21bai_2 _06868_ (.A1(_01137_),
    .A2(\rvsingle.dp.rf.rf[16][23] ),
    .B1_N(_01611_),
    .Y(_01789_));
 sky130_fd_sc_hd__and2b_2 _06869_ (.A_N(\rvsingle.dp.rf.rf[17][23] ),
    .B(_01558_),
    .X(_01790_));
 sky130_fd_sc_hd__o21ai_2 _06870_ (.A1(_01789_),
    .A2(_01790_),
    .B1(_01768_),
    .Y(_01791_));
 sky130_fd_sc_hd__or2b_2 _06871_ (.A(\rvsingle.dp.rf.rf[19][23] ),
    .B_N(_01753_),
    .X(_01792_));
 sky130_fd_sc_hd__o211a_2 _06872_ (.A1(_01126_),
    .A2(\rvsingle.dp.rf.rf[18][23] ),
    .B1(_01105_),
    .C1(_01792_),
    .X(_01793_));
 sky130_fd_sc_hd__nor2_2 _06873_ (.A(_01562_),
    .B(\rvsingle.dp.rf.rf[22][23] ),
    .Y(_01794_));
 sky130_fd_sc_hd__and2b_2 _06874_ (.A_N(\rvsingle.dp.rf.rf[23][23] ),
    .B(_01097_),
    .X(_01795_));
 sky130_fd_sc_hd__buf_1 _06875_ (.A(_01645_),
    .X(_01796_));
 sky130_fd_sc_hd__buf_1 _06876_ (.A(_01124_),
    .X(_01797_));
 sky130_fd_sc_hd__o21ba_2 _06877_ (.A1(_01797_),
    .A2(\rvsingle.dp.rf.rf[20][23] ),
    .B1_N(_01604_),
    .X(_01798_));
 sky130_fd_sc_hd__o21ai_2 _06878_ (.A1(_01796_),
    .A2(\rvsingle.dp.rf.rf[21][23] ),
    .B1(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__o311ai_2 _06879_ (.A1(_01668_),
    .A2(_01794_),
    .A3(_01795_),
    .B1(_01617_),
    .C1(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__o211ai_2 _06880_ (.A1(_01791_),
    .A2(_01793_),
    .B1(_01634_),
    .C1(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand3_2 _06881_ (.A(_01788_),
    .B(_01801_),
    .C(_01682_),
    .Y(_01802_));
 sky130_fd_sc_hd__nand4_2 _06882_ (.A(_01592_),
    .B(_01774_),
    .C(_01802_),
    .D(_01481_),
    .Y(_01803_));
 sky130_fd_sc_hd__and3_2 _06883_ (.A(_01591_),
    .B(_01580_),
    .C(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__mux4_2 _06884_ (.A0(\rvsingle.dp.rf.rf[12][23] ),
    .A1(\rvsingle.dp.rf.rf[13][23] ),
    .A2(\rvsingle.dp.rf.rf[14][23] ),
    .A3(\rvsingle.dp.rf.rf[15][23] ),
    .S0(_01417_),
    .S1(_01301_),
    .X(_01805_));
 sky130_fd_sc_hd__or2_2 _06885_ (.A(_01707_),
    .B(\rvsingle.dp.rf.rf[8][23] ),
    .X(_01806_));
 sky130_fd_sc_hd__o211ai_2 _06886_ (.A1(\rvsingle.dp.rf.rf[9][23] ),
    .A2(_01688_),
    .B1(_01689_),
    .C1(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__buf_1 _06887_ (.A(_01198_),
    .X(_01808_));
 sky130_fd_sc_hd__o21a_2 _06888_ (.A1(_01726_),
    .A2(\rvsingle.dp.rf.rf[10][23] ),
    .B1(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__o21ai_2 _06889_ (.A1(\rvsingle.dp.rf.rf[11][23] ),
    .A2(_01441_),
    .B1(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__a31oi_2 _06890_ (.A1(_01461_),
    .A2(_01807_),
    .A3(_01810_),
    .B1(_01218_),
    .Y(_01811_));
 sky130_fd_sc_hd__o21ai_2 _06891_ (.A1(_01208_),
    .A2(_01805_),
    .B1(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__mux4_2 _06892_ (.A0(\rvsingle.dp.rf.rf[0][23] ),
    .A1(\rvsingle.dp.rf.rf[1][23] ),
    .A2(\rvsingle.dp.rf.rf[2][23] ),
    .A3(\rvsingle.dp.rf.rf[3][23] ),
    .S0(_01469_),
    .S1(_01471_),
    .X(_01813_));
 sky130_fd_sc_hd__nor2_2 _06893_ (.A(_01336_),
    .B(\rvsingle.dp.rf.rf[4][23] ),
    .Y(_01814_));
 sky130_fd_sc_hd__o21ai_2 _06894_ (.A1(\rvsingle.dp.rf.rf[5][23] ),
    .A2(_01688_),
    .B1(_01689_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_2 _06895_ (.A(_01336_),
    .B(\rvsingle.dp.rf.rf[6][23] ),
    .Y(_01816_));
 sky130_fd_sc_hd__o21ai_2 _06896_ (.A1(\rvsingle.dp.rf.rf[7][23] ),
    .A2(_01688_),
    .B1(_01456_),
    .Y(_01817_));
 sky130_fd_sc_hd__o221ai_2 _06897_ (.A1(_01814_),
    .A2(_01815_),
    .B1(_01816_),
    .B2(_01817_),
    .C1(_01445_),
    .Y(_01818_));
 sky130_fd_sc_hd__o211ai_2 _06898_ (.A1(_01703_),
    .A2(_01813_),
    .B1(_01818_),
    .C1(_01218_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_2 _06899_ (.A(_01812_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__mux4_2 _06900_ (.A0(\rvsingle.dp.rf.rf[16][23] ),
    .A1(\rvsingle.dp.rf.rf[17][23] ),
    .A2(\rvsingle.dp.rf.rf[18][23] ),
    .A3(\rvsingle.dp.rf.rf[19][23] ),
    .S0(_01329_),
    .S1(_01456_),
    .X(_01821_));
 sky130_fd_sc_hd__nor2_2 _06901_ (.A(_01230_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__mux4_2 _06902_ (.A0(\rvsingle.dp.rf.rf[20][23] ),
    .A1(\rvsingle.dp.rf.rf[21][23] ),
    .A2(\rvsingle.dp.rf.rf[22][23] ),
    .A3(\rvsingle.dp.rf.rf[23][23] ),
    .S0(_01463_),
    .S1(_01471_),
    .X(_01823_));
 sky130_fd_sc_hd__o21ai_2 _06903_ (.A1(_01722_),
    .A2(_01823_),
    .B1(_01218_),
    .Y(_01824_));
 sky130_fd_sc_hd__mux4_2 _06904_ (.A0(\rvsingle.dp.rf.rf[28][23] ),
    .A1(\rvsingle.dp.rf.rf[29][23] ),
    .A2(\rvsingle.dp.rf.rf[30][23] ),
    .A3(\rvsingle.dp.rf.rf[31][23] ),
    .S0(_01463_),
    .S1(_01471_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_2 _06905_ (.A0(\rvsingle.dp.rf.rf[24][23] ),
    .A1(\rvsingle.dp.rf.rf[25][23] ),
    .S(_01335_),
    .X(_01826_));
 sky130_fd_sc_hd__buf_1 _06906_ (.A(_01294_),
    .X(_01827_));
 sky130_fd_sc_hd__buf_1 _06907_ (.A(_01190_),
    .X(_01828_));
 sky130_fd_sc_hd__or2_2 _06908_ (.A(_01828_),
    .B(\rvsingle.dp.rf.rf[26][23] ),
    .X(_01829_));
 sky130_fd_sc_hd__o211a_2 _06909_ (.A1(_01827_),
    .A2(\rvsingle.dp.rf.rf[27][23] ),
    .B1(_01808_),
    .C1(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__a211o_2 _06910_ (.A1(_01826_),
    .A2(_01309_),
    .B1(_01229_),
    .C1(_01830_),
    .X(_01831_));
 sky130_fd_sc_hd__o211ai_2 _06911_ (.A1(_01208_),
    .A2(_01825_),
    .B1(_01831_),
    .C1(_01478_),
    .Y(_01832_));
 sky130_fd_sc_hd__o211ai_2 _06912_ (.A1(_01822_),
    .A2(_01824_),
    .B1(_01188_),
    .C1(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__o211a_2 _06913_ (.A1(_01450_),
    .A2(_01820_),
    .B1(_01833_),
    .C1(_01247_),
    .X(_01834_));
 sky130_fd_sc_hd__a211o_2 _06914_ (.A1(_01587_),
    .A2(_01803_),
    .B1(_01066_),
    .C1(_01075_),
    .X(_01835_));
 sky130_fd_sc_hd__nand3b_2 _06915_ (.A_N(_01804_),
    .B(_01834_),
    .C(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__buf_1 _06916_ (.A(_01591_),
    .X(_01837_));
 sky130_fd_sc_hd__a21oi_2 _06917_ (.A1(_01581_),
    .A2(_01803_),
    .B1(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__o21bai_2 _06918_ (.A1(_01838_),
    .A2(_01804_),
    .B1_N(_01834_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_2 _06919_ (.A(_01836_),
    .B(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__nor2_2 _06920_ (.A(_01666_),
    .B(\rvsingle.dp.rf.rf[14][22] ),
    .Y(_01841_));
 sky130_fd_sc_hd__buf_1 _06921_ (.A(_01645_),
    .X(_01842_));
 sky130_fd_sc_hd__o21ai_2 _06922_ (.A1(\rvsingle.dp.rf.rf[15][22] ),
    .A2(_01842_),
    .B1(_01612_),
    .Y(_01843_));
 sky130_fd_sc_hd__nor2_2 _06923_ (.A(_01098_),
    .B(\rvsingle.dp.rf.rf[12][22] ),
    .Y(_01844_));
 sky130_fd_sc_hd__o21ai_2 _06924_ (.A1(\rvsingle.dp.rf.rf[13][22] ),
    .A2(_01088_),
    .B1(_01668_),
    .Y(_01845_));
 sky130_fd_sc_hd__o221a_2 _06925_ (.A1(_01841_),
    .A2(_01843_),
    .B1(_01844_),
    .B2(_01845_),
    .C1(_01112_),
    .X(_01846_));
 sky130_fd_sc_hd__buf_1 _06926_ (.A(_01752_),
    .X(_01847_));
 sky130_fd_sc_hd__buf_1 _06927_ (.A(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__or2b_2 _06928_ (.A(\rvsingle.dp.rf.rf[11][22] ),
    .B_N(_01097_),
    .X(_01849_));
 sky130_fd_sc_hd__o211ai_2 _06929_ (.A1(_01848_),
    .A2(\rvsingle.dp.rf.rf[10][22] ),
    .B1(_01612_),
    .C1(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__or2b_2 _06930_ (.A(\rvsingle.dp.rf.rf[9][22] ),
    .B_N(_01847_),
    .X(_01851_));
 sky130_fd_sc_hd__o211ai_2 _06931_ (.A1(_01848_),
    .A2(\rvsingle.dp.rf.rf[8][22] ),
    .B1(_01851_),
    .C1(_01759_),
    .Y(_01852_));
 sky130_fd_sc_hd__buf_1 _06932_ (.A(_01155_),
    .X(_01853_));
 sky130_fd_sc_hd__a31o_2 _06933_ (.A1(_01565_),
    .A2(_01850_),
    .A3(_01852_),
    .B1(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_2 _06934_ (.A0(\rvsingle.dp.rf.rf[0][22] ),
    .A1(\rvsingle.dp.rf.rf[1][22] ),
    .S(_01562_),
    .X(_01855_));
 sky130_fd_sc_hd__buf_1 _06935_ (.A(_01092_),
    .X(_01856_));
 sky130_fd_sc_hd__or2b_2 _06936_ (.A(\rvsingle.dp.rf.rf[3][22] ),
    .B_N(_01658_),
    .X(_01857_));
 sky130_fd_sc_hd__o211a_2 _06937_ (.A1(_01848_),
    .A2(\rvsingle.dp.rf.rf[2][22] ),
    .B1(_01612_),
    .C1(_01857_),
    .X(_01858_));
 sky130_fd_sc_hd__a211oi_2 _06938_ (.A1(_01855_),
    .A2(_01856_),
    .B1(_01512_),
    .C1(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__buf_1 _06939_ (.A(_01086_),
    .X(_01860_));
 sky130_fd_sc_hd__buf_1 _06940_ (.A(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__buf_1 _06941_ (.A(_01557_),
    .X(_01862_));
 sky130_fd_sc_hd__or2_2 _06942_ (.A(_01862_),
    .B(\rvsingle.dp.rf.rf[6][22] ),
    .X(_01863_));
 sky130_fd_sc_hd__o211ai_2 _06943_ (.A1(_01861_),
    .A2(\rvsingle.dp.rf.rf[7][22] ),
    .B1(_01655_),
    .C1(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__buf_1 _06944_ (.A(_01087_),
    .X(_01865_));
 sky130_fd_sc_hd__or2_2 _06945_ (.A(_01148_),
    .B(\rvsingle.dp.rf.rf[4][22] ),
    .X(_01866_));
 sky130_fd_sc_hd__o211ai_2 _06946_ (.A1(\rvsingle.dp.rf.rf[5][22] ),
    .A2(_01865_),
    .B1(_01759_),
    .C1(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__a31o_2 _06947_ (.A1(_01864_),
    .A2(_01867_),
    .A3(_01112_),
    .B1(_01116_),
    .X(_01868_));
 sky130_fd_sc_hd__o221ai_2 _06948_ (.A1(_01846_),
    .A2(_01854_),
    .B1(_01859_),
    .B2(_01868_),
    .C1(_01378_),
    .Y(_01869_));
 sky130_fd_sc_hd__buf_1 _06949_ (.A(_01082_),
    .X(_01870_));
 sky130_fd_sc_hd__nor2_2 _06950_ (.A(_01559_),
    .B(\rvsingle.dp.rf.rf[30][22] ),
    .Y(_01871_));
 sky130_fd_sc_hd__o21ai_2 _06951_ (.A1(\rvsingle.dp.rf.rf[31][22] ),
    .A2(_01865_),
    .B1(_01655_),
    .Y(_01872_));
 sky130_fd_sc_hd__or2_2 _06952_ (.A(_01862_),
    .B(\rvsingle.dp.rf.rf[28][22] ),
    .X(_01873_));
 sky130_fd_sc_hd__o211ai_2 _06953_ (.A1(\rvsingle.dp.rf.rf[29][22] ),
    .A2(_01861_),
    .B1(_01759_),
    .C1(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__o211a_2 _06954_ (.A1(_01871_),
    .A2(_01872_),
    .B1(_01112_),
    .C1(_01874_),
    .X(_01875_));
 sky130_fd_sc_hd__nor2_2 _06955_ (.A(_01744_),
    .B(\rvsingle.dp.rf.rf[24][22] ),
    .Y(_01876_));
 sky130_fd_sc_hd__buf_1 _06956_ (.A(_01095_),
    .X(_01877_));
 sky130_fd_sc_hd__buf_1 _06957_ (.A(_01877_),
    .X(_01878_));
 sky130_fd_sc_hd__and2b_2 _06958_ (.A_N(\rvsingle.dp.rf.rf[25][22] ),
    .B(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__buf_1 _06959_ (.A(_01258_),
    .X(_01880_));
 sky130_fd_sc_hd__o21a_2 _06960_ (.A1(_01558_),
    .A2(\rvsingle.dp.rf.rf[26][22] ),
    .B1(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__o21ai_2 _06961_ (.A1(\rvsingle.dp.rf.rf[27][22] ),
    .A2(_01865_),
    .B1(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__o311ai_2 _06962_ (.A1(_01260_),
    .A2(_01876_),
    .A3(_01879_),
    .B1(_01565_),
    .C1(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__nand2_2 _06963_ (.A(_01883_),
    .B(_01526_),
    .Y(_01884_));
 sky130_fd_sc_hd__nor2_2 _06964_ (.A(_01098_),
    .B(\rvsingle.dp.rf.rf[18][22] ),
    .Y(_01885_));
 sky130_fd_sc_hd__o21ai_2 _06965_ (.A1(\rvsingle.dp.rf.rf[19][22] ),
    .A2(_01088_),
    .B1(_01626_),
    .Y(_01886_));
 sky130_fd_sc_hd__or2_2 _06966_ (.A(_01642_),
    .B(\rvsingle.dp.rf.rf[16][22] ),
    .X(_01887_));
 sky130_fd_sc_hd__o211ai_2 _06967_ (.A1(\rvsingle.dp.rf.rf[17][22] ),
    .A2(_01088_),
    .B1(_01092_),
    .C1(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__o211ai_2 _06968_ (.A1(_01885_),
    .A2(_01886_),
    .B1(_01888_),
    .C1(_01565_),
    .Y(_01889_));
 sky130_fd_sc_hd__nor2_2 _06969_ (.A(_01098_),
    .B(\rvsingle.dp.rf.rf[22][22] ),
    .Y(_01890_));
 sky130_fd_sc_hd__o21ai_2 _06970_ (.A1(\rvsingle.dp.rf.rf[23][22] ),
    .A2(_01865_),
    .B1(_01626_),
    .Y(_01891_));
 sky130_fd_sc_hd__or2_2 _06971_ (.A(_01675_),
    .B(\rvsingle.dp.rf.rf[20][22] ),
    .X(_01892_));
 sky130_fd_sc_hd__o211ai_2 _06972_ (.A1(\rvsingle.dp.rf.rf[21][22] ),
    .A2(_01865_),
    .B1(_01668_),
    .C1(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__o211ai_2 _06973_ (.A1(_01890_),
    .A2(_01891_),
    .B1(_01503_),
    .C1(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand3_2 _06974_ (.A(_01157_),
    .B(_01889_),
    .C(_01894_),
    .Y(_01895_));
 sky130_fd_sc_hd__o211ai_2 _06975_ (.A1(_01875_),
    .A2(_01884_),
    .B1(_01682_),
    .C1(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__nand4_2 _06976_ (.A(_01869_),
    .B(_01870_),
    .C(_01592_),
    .D(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__and3_2 _06977_ (.A(_01591_),
    .B(_01580_),
    .C(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__mux4_2 _06978_ (.A0(\rvsingle.dp.rf.rf[20][22] ),
    .A1(\rvsingle.dp.rf.rf[21][22] ),
    .A2(\rvsingle.dp.rf.rf[22][22] ),
    .A3(\rvsingle.dp.rf.rf[23][22] ),
    .S0(_01417_),
    .S1(_01301_),
    .X(_01899_));
 sky130_fd_sc_hd__nor2_2 _06979_ (.A(_01329_),
    .B(\rvsingle.dp.rf.rf[18][22] ),
    .Y(_01900_));
 sky130_fd_sc_hd__buf_1 _06980_ (.A(_01294_),
    .X(_01901_));
 sky130_fd_sc_hd__o21ai_2 _06981_ (.A1(\rvsingle.dp.rf.rf[19][22] ),
    .A2(_01901_),
    .B1(_01244_),
    .Y(_01902_));
 sky130_fd_sc_hd__buf_1 _06982_ (.A(_01327_),
    .X(_01903_));
 sky130_fd_sc_hd__or2_2 _06983_ (.A(_01903_),
    .B(\rvsingle.dp.rf.rf[16][22] ),
    .X(_01904_));
 sky130_fd_sc_hd__o211ai_2 _06984_ (.A1(\rvsingle.dp.rf.rf[17][22] ),
    .A2(_01424_),
    .B1(_01716_),
    .C1(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__o211a_2 _06985_ (.A1(_01900_),
    .A2(_01902_),
    .B1(_01721_),
    .C1(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__o21bai_2 _06986_ (.A1(_01208_),
    .A2(_01899_),
    .B1_N(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__mux4_2 _06987_ (.A0(\rvsingle.dp.rf.rf[28][22] ),
    .A1(\rvsingle.dp.rf.rf[29][22] ),
    .A2(\rvsingle.dp.rf.rf[30][22] ),
    .A3(\rvsingle.dp.rf.rf[31][22] ),
    .S0(_01329_),
    .S1(_01456_),
    .X(_01908_));
 sky130_fd_sc_hd__or2_2 _06988_ (.A(_01469_),
    .B(\rvsingle.dp.rf.rf[26][22] ),
    .X(_01909_));
 sky130_fd_sc_hd__o211a_2 _06989_ (.A1(_01296_),
    .A2(\rvsingle.dp.rf.rf[27][22] ),
    .B1(_01434_),
    .C1(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_2 _06990_ (.A0(\rvsingle.dp.rf.rf[24][22] ),
    .A1(\rvsingle.dp.rf.rf[25][22] ),
    .S(_01695_),
    .X(_01911_));
 sky130_fd_sc_hd__a21o_2 _06991_ (.A1(_01911_),
    .A2(_01309_),
    .B1(_01711_),
    .X(_01912_));
 sky130_fd_sc_hd__o221ai_2 _06992_ (.A1(_01208_),
    .A2(_01908_),
    .B1(_01910_),
    .B2(_01912_),
    .C1(_01222_),
    .Y(_01913_));
 sky130_fd_sc_hd__o21ai_2 _06993_ (.A1(_01222_),
    .A2(_01907_),
    .B1(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__buf_1 _06994_ (.A(_01694_),
    .X(_01915_));
 sky130_fd_sc_hd__mux4_2 _06995_ (.A0(\rvsingle.dp.rf.rf[8][22] ),
    .A1(\rvsingle.dp.rf.rf[9][22] ),
    .A2(\rvsingle.dp.rf.rf[10][22] ),
    .A3(\rvsingle.dp.rf.rf[11][22] ),
    .S0(_01242_),
    .S1(_01434_),
    .X(_01916_));
 sky130_fd_sc_hd__mux4_2 _06996_ (.A0(\rvsingle.dp.rf.rf[12][22] ),
    .A1(\rvsingle.dp.rf.rf[13][22] ),
    .A2(\rvsingle.dp.rf.rf[14][22] ),
    .A3(\rvsingle.dp.rf.rf[15][22] ),
    .S0(_01335_),
    .S1(_01199_),
    .X(_01917_));
 sky130_fd_sc_hd__o21a_2 _06997_ (.A1(_01461_),
    .A2(_01917_),
    .B1(_01447_),
    .X(_01918_));
 sky130_fd_sc_hd__o21ai_2 _06998_ (.A1(_01915_),
    .A2(_01916_),
    .B1(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__mux4_2 _06999_ (.A0(\rvsingle.dp.rf.rf[0][22] ),
    .A1(\rvsingle.dp.rf.rf[1][22] ),
    .A2(\rvsingle.dp.rf.rf[2][22] ),
    .A3(\rvsingle.dp.rf.rf[3][22] ),
    .S0(_01432_),
    .S1(_01434_),
    .X(_01920_));
 sky130_fd_sc_hd__mux4_2 _07000_ (.A0(\rvsingle.dp.rf.rf[4][22] ),
    .A1(\rvsingle.dp.rf.rf[5][22] ),
    .A2(\rvsingle.dp.rf.rf[6][22] ),
    .A3(\rvsingle.dp.rf.rf[7][22] ),
    .S0(_01335_),
    .S1(_01199_),
    .X(_01921_));
 sky130_fd_sc_hd__o21a_2 _07001_ (.A1(_01461_),
    .A2(_01921_),
    .B1(_01699_),
    .X(_01922_));
 sky130_fd_sc_hd__o21ai_2 _07002_ (.A1(_01915_),
    .A2(_01920_),
    .B1(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__nand3_2 _07003_ (.A(_01316_),
    .B(_01919_),
    .C(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__o211a_2 _07004_ (.A1(_01317_),
    .A2(_01914_),
    .B1(_01924_),
    .C1(_01247_),
    .X(_01925_));
 sky130_fd_sc_hd__a211o_2 _07005_ (.A1(_01587_),
    .A2(_01897_),
    .B1(_01066_),
    .C1(_01075_),
    .X(_01926_));
 sky130_fd_sc_hd__nand3b_2 _07006_ (.A_N(_01898_),
    .B(_01925_),
    .C(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__a21oi_2 _07007_ (.A1(_01581_),
    .A2(_01897_),
    .B1(_01837_),
    .Y(_01928_));
 sky130_fd_sc_hd__o21bai_2 _07008_ (.A1(_01928_),
    .A2(_01898_),
    .B1_N(_01925_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_2 _07009_ (.A(_01927_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__nor4_2 _07010_ (.A(_01590_),
    .B(_01742_),
    .C(_01840_),
    .D(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__mux4_2 _07011_ (.A0(\rvsingle.dp.rf.rf[20][19] ),
    .A1(\rvsingle.dp.rf.rf[21][19] ),
    .A2(\rvsingle.dp.rf.rf[22][19] ),
    .A3(\rvsingle.dp.rf.rf[23][19] ),
    .S0(_01463_),
    .S1(_01456_),
    .X(_01932_));
 sky130_fd_sc_hd__nor2_2 _07012_ (.A(_01722_),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__mux4_2 _07013_ (.A0(\rvsingle.dp.rf.rf[16][19] ),
    .A1(\rvsingle.dp.rf.rf[17][19] ),
    .A2(\rvsingle.dp.rf.rf[18][19] ),
    .A3(\rvsingle.dp.rf.rf[19][19] ),
    .S0(_01329_),
    .S1(_01456_),
    .X(_01934_));
 sky130_fd_sc_hd__nor2_2 _07014_ (.A(_01230_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__mux4_2 _07015_ (.A0(\rvsingle.dp.rf.rf[24][19] ),
    .A1(\rvsingle.dp.rf.rf[25][19] ),
    .A2(\rvsingle.dp.rf.rf[26][19] ),
    .A3(\rvsingle.dp.rf.rf[27][19] ),
    .S0(_01469_),
    .S1(_01728_),
    .X(_01936_));
 sky130_fd_sc_hd__or2_2 _07016_ (.A(_01695_),
    .B(\rvsingle.dp.rf.rf[30][19] ),
    .X(_01937_));
 sky130_fd_sc_hd__o211a_2 _07017_ (.A1(_01441_),
    .A2(\rvsingle.dp.rf.rf[31][19] ),
    .B1(_01301_),
    .C1(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_2 _07018_ (.A0(\rvsingle.dp.rf.rf[28][19] ),
    .A1(\rvsingle.dp.rf.rf[29][19] ),
    .S(_01691_),
    .X(_01939_));
 sky130_fd_sc_hd__a21o_2 _07019_ (.A1(_01939_),
    .A2(_01309_),
    .B1(_01207_),
    .X(_01940_));
 sky130_fd_sc_hd__o221ai_2 _07020_ (.A1(_01703_),
    .A2(_01936_),
    .B1(_01938_),
    .B2(_01940_),
    .C1(_01478_),
    .Y(_01941_));
 sky130_fd_sc_hd__o311ai_2 _07021_ (.A1(_01222_),
    .A2(_01933_),
    .A3(_01935_),
    .B1(_01450_),
    .C1(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__buf_1 _07022_ (.A(_01424_),
    .X(_01943_));
 sky130_fd_sc_hd__o21a_2 _07023_ (.A1(_01242_),
    .A2(\rvsingle.dp.rf.rf[10][19] ),
    .B1(_01728_),
    .X(_01944_));
 sky130_fd_sc_hd__o21ai_2 _07024_ (.A1(\rvsingle.dp.rf.rf[11][19] ),
    .A2(_01943_),
    .B1(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__mux2_2 _07025_ (.A0(\rvsingle.dp.rf.rf[8][19] ),
    .A1(\rvsingle.dp.rf.rf[9][19] ),
    .S(_01469_),
    .X(_01946_));
 sky130_fd_sc_hd__a21oi_2 _07026_ (.A1(_01946_),
    .A2(_01717_),
    .B1(_01445_),
    .Y(_01947_));
 sky130_fd_sc_hd__mux4_2 _07027_ (.A0(\rvsingle.dp.rf.rf[12][19] ),
    .A1(\rvsingle.dp.rf.rf[13][19] ),
    .A2(\rvsingle.dp.rf.rf[14][19] ),
    .A3(\rvsingle.dp.rf.rf[15][19] ),
    .S0(_01329_),
    .S1(_01456_),
    .X(_01948_));
 sky130_fd_sc_hd__o2bb2ai_2 _07028_ (.A1_N(_01945_),
    .A2_N(_01947_),
    .B1(_01208_),
    .B2(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__mux4_2 _07029_ (.A0(\rvsingle.dp.rf.rf[4][19] ),
    .A1(\rvsingle.dp.rf.rf[5][19] ),
    .A2(\rvsingle.dp.rf.rf[6][19] ),
    .A3(\rvsingle.dp.rf.rf[7][19] ),
    .S0(_01417_),
    .S1(_01301_),
    .X(_01950_));
 sky130_fd_sc_hd__or2_2 _07030_ (.A(_01707_),
    .B(\rvsingle.dp.rf.rf[0][19] ),
    .X(_01951_));
 sky130_fd_sc_hd__o211ai_2 _07031_ (.A1(\rvsingle.dp.rf.rf[1][19] ),
    .A2(_01441_),
    .B1(_01689_),
    .C1(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__buf_1 _07032_ (.A(_01198_),
    .X(_01953_));
 sky130_fd_sc_hd__o21a_2 _07033_ (.A1(_01726_),
    .A2(\rvsingle.dp.rf.rf[2][19] ),
    .B1(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__o21ai_2 _07034_ (.A1(\rvsingle.dp.rf.rf[3][19] ),
    .A2(_01441_),
    .B1(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__a31oi_2 _07035_ (.A1(_01461_),
    .A2(_01952_),
    .A3(_01955_),
    .B1(_01447_),
    .Y(_01956_));
 sky130_fd_sc_hd__o21ai_2 _07036_ (.A1(_01208_),
    .A2(_01950_),
    .B1(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__o211ai_2 _07037_ (.A1(_01218_),
    .A2(_01949_),
    .B1(_01957_),
    .C1(_01316_),
    .Y(_01958_));
 sky130_fd_sc_hd__and3_2 _07038_ (.A(_01247_),
    .B(_01942_),
    .C(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__buf_1 _07039_ (.A(_01064_),
    .X(_01960_));
 sky130_fd_sc_hd__buf_1 _07040_ (.A(_01177_),
    .X(_01961_));
 sky130_fd_sc_hd__buf_1 _07041_ (.A(_01150_),
    .X(_01962_));
 sky130_fd_sc_hd__nor2_2 _07042_ (.A(_01656_),
    .B(\rvsingle.dp.rf.rf[16][19] ),
    .Y(_01963_));
 sky130_fd_sc_hd__and2b_2 _07043_ (.A_N(\rvsingle.dp.rf.rf[17][19] ),
    .B(_01862_),
    .X(_01964_));
 sky130_fd_sc_hd__or2b_2 _07044_ (.A(\rvsingle.dp.rf.rf[19][19] ),
    .B_N(_01650_),
    .X(_01965_));
 sky130_fd_sc_hd__o211ai_2 _07045_ (.A1(_01256_),
    .A2(\rvsingle.dp.rf.rf[18][19] ),
    .B1(_01660_),
    .C1(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__o311ai_2 _07046_ (.A1(_01655_),
    .A2(_01963_),
    .A3(_01964_),
    .B1(_01768_),
    .C1(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__o21ba_2 _07047_ (.A1(_01658_),
    .A2(\rvsingle.dp.rf.rf[20][19] ),
    .B1_N(_01647_),
    .X(_01968_));
 sky130_fd_sc_hd__o21ai_2 _07048_ (.A1(_01088_),
    .A2(\rvsingle.dp.rf.rf[21][19] ),
    .B1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__o21a_2 _07049_ (.A1(_01148_),
    .A2(\rvsingle.dp.rf.rf[22][19] ),
    .B1(_01611_),
    .X(_01970_));
 sky130_fd_sc_hd__o21ai_2 _07050_ (.A1(\rvsingle.dp.rf.rf[23][19] ),
    .A2(_01842_),
    .B1(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__nand3_2 _07051_ (.A(_01969_),
    .B(_01632_),
    .C(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__nand3_2 _07052_ (.A(_01634_),
    .B(_01967_),
    .C(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor2_2 _07053_ (.A(_01656_),
    .B(\rvsingle.dp.rf.rf[24][19] ),
    .Y(_01974_));
 sky130_fd_sc_hd__and2b_2 _07054_ (.A_N(\rvsingle.dp.rf.rf[25][19] ),
    .B(_01862_),
    .X(_01975_));
 sky130_fd_sc_hd__or2b_2 _07055_ (.A(\rvsingle.dp.rf.rf[27][19] ),
    .B_N(_01650_),
    .X(_01976_));
 sky130_fd_sc_hd__o211ai_2 _07056_ (.A1(_01256_),
    .A2(\rvsingle.dp.rf.rf[26][19] ),
    .B1(_01660_),
    .C1(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__o311ai_2 _07057_ (.A1(_01655_),
    .A2(_01974_),
    .A3(_01975_),
    .B1(_01768_),
    .C1(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__o21ba_2 _07058_ (.A1(_01675_),
    .A2(\rvsingle.dp.rf.rf[28][19] ),
    .B1_N(_01104_),
    .X(_01979_));
 sky130_fd_sc_hd__o21ai_2 _07059_ (.A1(_01842_),
    .A2(\rvsingle.dp.rf.rf[29][19] ),
    .B1(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__o21a_2 _07060_ (.A1(_01642_),
    .A2(\rvsingle.dp.rf.rf[30][19] ),
    .B1(_01596_),
    .X(_01981_));
 sky130_fd_sc_hd__o21ai_2 _07061_ (.A1(\rvsingle.dp.rf.rf[31][19] ),
    .A2(_01842_),
    .B1(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand3_2 _07062_ (.A(_01980_),
    .B(_01632_),
    .C(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand3_2 _07063_ (.A(_01978_),
    .B(_01983_),
    .C(_01116_),
    .Y(_01984_));
 sky130_fd_sc_hd__nand3_2 _07064_ (.A(_01973_),
    .B(_01682_),
    .C(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__nor2_2 _07065_ (.A(_01603_),
    .B(\rvsingle.dp.rf.rf[8][19] ),
    .Y(_01986_));
 sky130_fd_sc_hd__and2b_2 _07066_ (.A_N(\rvsingle.dp.rf.rf[9][19] ),
    .B(_01382_),
    .X(_01987_));
 sky130_fd_sc_hd__or2b_2 _07067_ (.A(\rvsingle.dp.rf.rf[11][19] ),
    .B_N(_01753_),
    .X(_01988_));
 sky130_fd_sc_hd__o211ai_2 _07068_ (.A1(_01744_),
    .A2(\rvsingle.dp.rf.rf[10][19] ),
    .B1(_01648_),
    .C1(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__o311a_2 _07069_ (.A1(_01655_),
    .A2(_01986_),
    .A3(_01987_),
    .B1(_01768_),
    .C1(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__inv_2 _07070_ (.A(\rvsingle.dp.rf.rf[15][19] ),
    .Y(_01991_));
 sky130_fd_sc_hd__o21ai_2 _07071_ (.A1(_01656_),
    .A2(\rvsingle.dp.rf.rf[14][19] ),
    .B1(_01605_),
    .Y(_01992_));
 sky130_fd_sc_hd__a21oi_2 _07072_ (.A1(_01991_),
    .A2(_01383_),
    .B1(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__o21bai_2 _07073_ (.A1(_01518_),
    .A2(\rvsingle.dp.rf.rf[12][19] ),
    .B1_N(_01611_),
    .Y(_01994_));
 sky130_fd_sc_hd__and2b_2 _07074_ (.A_N(\rvsingle.dp.rf.rf[13][19] ),
    .B(_01630_),
    .X(_01995_));
 sky130_fd_sc_hd__o21ai_2 _07075_ (.A1(_01994_),
    .A2(_01995_),
    .B1(_01632_),
    .Y(_01996_));
 sky130_fd_sc_hd__o21ai_2 _07076_ (.A1(_01993_),
    .A2(_01996_),
    .B1(_01116_),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_2 _07077_ (.A(_01614_),
    .B(\rvsingle.dp.rf.rf[0][19] ),
    .Y(_01998_));
 sky130_fd_sc_hd__and2b_2 _07078_ (.A_N(\rvsingle.dp.rf.rf[1][19] ),
    .B(_01847_),
    .X(_01999_));
 sky130_fd_sc_hd__or2b_2 _07079_ (.A(\rvsingle.dp.rf.rf[3][19] ),
    .B_N(_01255_),
    .X(_02000_));
 sky130_fd_sc_hd__o211ai_2 _07080_ (.A1(_01619_),
    .A2(\rvsingle.dp.rf.rf[2][19] ),
    .B1(_01620_),
    .C1(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__o311ai_2 _07081_ (.A1(_01648_),
    .A2(_01998_),
    .A3(_01999_),
    .B1(_01600_),
    .C1(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__nor2_2 _07082_ (.A(_01614_),
    .B(\rvsingle.dp.rf.rf[6][19] ),
    .Y(_02003_));
 sky130_fd_sc_hd__and2b_2 _07083_ (.A_N(\rvsingle.dp.rf.rf[7][19] ),
    .B(_01675_),
    .X(_02004_));
 sky130_fd_sc_hd__buf_1 _07084_ (.A(_01124_),
    .X(_02005_));
 sky130_fd_sc_hd__o21ba_2 _07085_ (.A1(_02005_),
    .A2(\rvsingle.dp.rf.rf[4][19] ),
    .B1_N(_01530_),
    .X(_02006_));
 sky130_fd_sc_hd__o21ai_2 _07086_ (.A1(_01796_),
    .A2(\rvsingle.dp.rf.rf[5][19] ),
    .B1(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__o311ai_2 _07087_ (.A1(_01092_),
    .A2(_02003_),
    .A3(_02004_),
    .B1(_01617_),
    .C1(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand3_2 _07088_ (.A(_01634_),
    .B(_02002_),
    .C(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__o211ai_2 _07089_ (.A1(_01990_),
    .A2(_01997_),
    .B1(_02009_),
    .C1(_01593_),
    .Y(_02010_));
 sky130_fd_sc_hd__o211ai_2 _07090_ (.A1(_01962_),
    .A2(_01128_),
    .B1(_01985_),
    .C1(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__o221ai_2 _07091_ (.A1(_01960_),
    .A2(_01075_),
    .B1(_01961_),
    .B2(_02011_),
    .C1(_01587_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand2_2 _07092_ (.A(_02011_),
    .B(_01084_),
    .Y(_02013_));
 sky130_fd_sc_hd__o211ai_2 _07093_ (.A1(_01482_),
    .A2(_01171_),
    .B1(_01584_),
    .C1(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__nand3_2 _07094_ (.A(_01959_),
    .B(_02012_),
    .C(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__a32o_2 _07095_ (.A1(_01248_),
    .A2(_01942_),
    .A3(_01958_),
    .B1(_02012_),
    .B2(_02014_),
    .X(_02016_));
 sky130_fd_sc_hd__nor2_2 _07096_ (.A(_01383_),
    .B(\rvsingle.dp.rf.rf[24][18] ),
    .Y(_02017_));
 sky130_fd_sc_hd__o21ai_2 _07097_ (.A1(\rvsingle.dp.rf.rf[25][18] ),
    .A2(_01861_),
    .B1(_01759_),
    .Y(_02018_));
 sky130_fd_sc_hd__o21a_2 _07098_ (.A1(_01595_),
    .A2(\rvsingle.dp.rf.rf[26][18] ),
    .B1(_01490_),
    .X(_02019_));
 sky130_fd_sc_hd__o21ai_2 _07099_ (.A1(\rvsingle.dp.rf.rf[27][18] ),
    .A2(_01540_),
    .B1(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__o211ai_2 _07100_ (.A1(_02017_),
    .A2(_02018_),
    .B1(_01132_),
    .C1(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__nor2_2 _07101_ (.A(_01559_),
    .B(\rvsingle.dp.rf.rf[30][18] ),
    .Y(_02022_));
 sky130_fd_sc_hd__o21ai_2 _07102_ (.A1(\rvsingle.dp.rf.rf[31][18] ),
    .A2(_01865_),
    .B1(_01655_),
    .Y(_02023_));
 sky130_fd_sc_hd__or2_2 _07103_ (.A(_01097_),
    .B(\rvsingle.dp.rf.rf[28][18] ),
    .X(_02024_));
 sky130_fd_sc_hd__o211ai_2 _07104_ (.A1(\rvsingle.dp.rf.rf[29][18] ),
    .A2(_01861_),
    .B1(_01759_),
    .C1(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__o211ai_2 _07105_ (.A1(_02022_),
    .A2(_02023_),
    .B1(_01112_),
    .C1(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__nand3_2 _07106_ (.A(_02021_),
    .B(_02026_),
    .C(_01526_),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_2 _07107_ (.A(_01666_),
    .B(\rvsingle.dp.rf.rf[16][18] ),
    .Y(_02028_));
 sky130_fd_sc_hd__o21ai_2 _07108_ (.A1(\rvsingle.dp.rf.rf[17][18] ),
    .A2(_01088_),
    .B1(_01668_),
    .Y(_02029_));
 sky130_fd_sc_hd__buf_1 _07109_ (.A(_01566_),
    .X(_02030_));
 sky130_fd_sc_hd__buf_1 _07110_ (.A(_01258_),
    .X(_02031_));
 sky130_fd_sc_hd__o21a_2 _07111_ (.A1(_02030_),
    .A2(\rvsingle.dp.rf.rf[18][18] ),
    .B1(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__o21ai_2 _07112_ (.A1(\rvsingle.dp.rf.rf[19][18] ),
    .A2(_01861_),
    .B1(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__o211ai_2 _07113_ (.A1(_02028_),
    .A2(_02029_),
    .B1(_01565_),
    .C1(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__nor2_2 _07114_ (.A(_01744_),
    .B(\rvsingle.dp.rf.rf[20][18] ),
    .Y(_02035_));
 sky130_fd_sc_hd__and2b_2 _07115_ (.A_N(\rvsingle.dp.rf.rf[21][18] ),
    .B(_01878_),
    .X(_02036_));
 sky130_fd_sc_hd__o21a_2 _07116_ (.A1(_01558_),
    .A2(\rvsingle.dp.rf.rf[22][18] ),
    .B1(_01880_),
    .X(_02037_));
 sky130_fd_sc_hd__o21ai_2 _07117_ (.A1(\rvsingle.dp.rf.rf[23][18] ),
    .A2(_01865_),
    .B1(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__o311ai_2 _07118_ (.A1(_01260_),
    .A2(_02035_),
    .A3(_02036_),
    .B1(_01503_),
    .C1(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand3_2 _07119_ (.A(_01634_),
    .B(_02034_),
    .C(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__nand3_2 _07120_ (.A(_02027_),
    .B(_02040_),
    .C(_01682_),
    .Y(_02041_));
 sky130_fd_sc_hd__nor2_2 _07121_ (.A(_01383_),
    .B(\rvsingle.dp.rf.rf[6][18] ),
    .Y(_02042_));
 sky130_fd_sc_hd__o21ai_2 _07122_ (.A1(\rvsingle.dp.rf.rf[7][18] ),
    .A2(_01861_),
    .B1(_01260_),
    .Y(_02043_));
 sky130_fd_sc_hd__or2_2 _07123_ (.A(_01630_),
    .B(\rvsingle.dp.rf.rf[4][18] ),
    .X(_02044_));
 sky130_fd_sc_hd__o211ai_2 _07124_ (.A1(\rvsingle.dp.rf.rf[5][18] ),
    .A2(_01540_),
    .B1(_01759_),
    .C1(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__o211a_2 _07125_ (.A1(_02042_),
    .A2(_02043_),
    .B1(_02045_),
    .C1(_01112_),
    .X(_02046_));
 sky130_fd_sc_hd__or2b_2 _07126_ (.A(\rvsingle.dp.rf.rf[3][18] ),
    .B_N(_01567_),
    .X(_02047_));
 sky130_fd_sc_hd__o211ai_2 _07127_ (.A1(_01559_),
    .A2(\rvsingle.dp.rf.rf[2][18] ),
    .B1(_01260_),
    .C1(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__or2b_2 _07128_ (.A(\rvsingle.dp.rf.rf[1][18] ),
    .B_N(_01558_),
    .X(_02049_));
 sky130_fd_sc_hd__o211ai_2 _07129_ (.A1(_01559_),
    .A2(\rvsingle.dp.rf.rf[0][18] ),
    .B1(_02049_),
    .C1(_01543_),
    .Y(_02050_));
 sky130_fd_sc_hd__a31o_2 _07130_ (.A1(_01132_),
    .A2(_02048_),
    .A3(_02050_),
    .B1(_01116_),
    .X(_02051_));
 sky130_fd_sc_hd__nor2_2 _07131_ (.A(_01383_),
    .B(\rvsingle.dp.rf.rf[12][18] ),
    .Y(_02052_));
 sky130_fd_sc_hd__o21ai_2 _07132_ (.A1(\rvsingle.dp.rf.rf[13][18] ),
    .A2(_01540_),
    .B1(_01543_),
    .Y(_02053_));
 sky130_fd_sc_hd__o21a_2 _07133_ (.A1(_01493_),
    .A2(\rvsingle.dp.rf.rf[14][18] ),
    .B1(_01523_),
    .X(_02054_));
 sky130_fd_sc_hd__o21ai_2 _07134_ (.A1(\rvsingle.dp.rf.rf[15][18] ),
    .A2(_01509_),
    .B1(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__o211ai_2 _07135_ (.A1(_02052_),
    .A2(_02053_),
    .B1(_01112_),
    .C1(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_2 _07136_ (.A(_01559_),
    .B(\rvsingle.dp.rf.rf[8][18] ),
    .Y(_02057_));
 sky130_fd_sc_hd__o21ai_2 _07137_ (.A1(\rvsingle.dp.rf.rf[9][18] ),
    .A2(_01861_),
    .B1(_01759_),
    .Y(_02058_));
 sky130_fd_sc_hd__buf_1 _07138_ (.A(_01519_),
    .X(_02059_));
 sky130_fd_sc_hd__o21a_2 _07139_ (.A1(_01268_),
    .A2(\rvsingle.dp.rf.rf[10][18] ),
    .B1(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__o21ai_2 _07140_ (.A1(\rvsingle.dp.rf.rf[11][18] ),
    .A2(_01540_),
    .B1(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__o211ai_2 _07141_ (.A1(_02057_),
    .A2(_02058_),
    .B1(_01565_),
    .C1(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand3_2 _07142_ (.A(_02056_),
    .B(_02062_),
    .C(_01506_),
    .Y(_02063_));
 sky130_fd_sc_hd__o211ai_2 _07143_ (.A1(_02046_),
    .A2(_02051_),
    .B1(_01593_),
    .C1(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__o211ai_2 _07144_ (.A1(_01962_),
    .A2(_01100_),
    .B1(_02041_),
    .C1(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__o221ai_2 _07145_ (.A1(_01960_),
    .A2(_01075_),
    .B1(_01961_),
    .B2(_02065_),
    .C1(_01587_),
    .Y(_02066_));
 sky130_fd_sc_hd__nand4_2 _07146_ (.A(_02064_),
    .B(_01870_),
    .C(_01153_),
    .D(_02041_),
    .Y(_02067_));
 sky130_fd_sc_hd__a21o_2 _07147_ (.A1(_01587_),
    .A2(_02067_),
    .B1(_01486_),
    .X(_02068_));
 sky130_fd_sc_hd__mux4_2 _07148_ (.A0(\rvsingle.dp.rf.rf[0][18] ),
    .A1(\rvsingle.dp.rf.rf[1][18] ),
    .A2(\rvsingle.dp.rf.rf[2][18] ),
    .A3(\rvsingle.dp.rf.rf[3][18] ),
    .S0(_01193_),
    .S1(_01451_),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_2 _07149_ (.A0(\rvsingle.dp.rf.rf[4][18] ),
    .A1(\rvsingle.dp.rf.rf[5][18] ),
    .S(_01432_),
    .X(_02070_));
 sky130_fd_sc_hd__or2_2 _07150_ (.A(_01695_),
    .B(\rvsingle.dp.rf.rf[6][18] ),
    .X(_02071_));
 sky130_fd_sc_hd__o211a_2 _07151_ (.A1(_01688_),
    .A2(\rvsingle.dp.rf.rf[7][18] ),
    .B1(_01301_),
    .C1(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__a211o_2 _07152_ (.A1(_02070_),
    .A2(_01717_),
    .B1(_01722_),
    .C1(_02072_),
    .X(_02073_));
 sky130_fd_sc_hd__o21ai_2 _07153_ (.A1(_01915_),
    .A2(_02069_),
    .B1(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__mux4_2 _07154_ (.A0(\rvsingle.dp.rf.rf[8][18] ),
    .A1(\rvsingle.dp.rf.rf[9][18] ),
    .A2(\rvsingle.dp.rf.rf[10][18] ),
    .A3(\rvsingle.dp.rf.rf[11][18] ),
    .S0(_01336_),
    .S1(_01200_),
    .X(_02075_));
 sky130_fd_sc_hd__or2_2 _07155_ (.A(_01336_),
    .B(\rvsingle.dp.rf.rf[14][18] ),
    .X(_02076_));
 sky130_fd_sc_hd__o211a_2 _07156_ (.A1(_01943_),
    .A2(\rvsingle.dp.rf.rf[15][18] ),
    .B1(_01451_),
    .C1(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_2 _07157_ (.A0(\rvsingle.dp.rf.rf[12][18] ),
    .A1(\rvsingle.dp.rf.rf[13][18] ),
    .S(_01432_),
    .X(_02078_));
 sky130_fd_sc_hd__a21o_2 _07158_ (.A1(_02078_),
    .A2(_01717_),
    .B1(_01722_),
    .X(_02079_));
 sky130_fd_sc_hd__o221ai_2 _07159_ (.A1(_01915_),
    .A2(_02075_),
    .B1(_02077_),
    .B2(_02079_),
    .C1(_01222_),
    .Y(_02080_));
 sky130_fd_sc_hd__o211a_2 _07160_ (.A1(_01223_),
    .A2(_02074_),
    .B1(_02080_),
    .C1(_01317_),
    .X(_02081_));
 sky130_fd_sc_hd__mux4_2 _07161_ (.A0(\rvsingle.dp.rf.rf[16][18] ),
    .A1(\rvsingle.dp.rf.rf[17][18] ),
    .A2(\rvsingle.dp.rf.rf[18][18] ),
    .A3(\rvsingle.dp.rf.rf[19][18] ),
    .S0(_01242_),
    .S1(_01434_),
    .X(_02082_));
 sky130_fd_sc_hd__nor2_2 _07162_ (.A(_01330_),
    .B(\rvsingle.dp.rf.rf[20][18] ),
    .Y(_02083_));
 sky130_fd_sc_hd__o21ai_2 _07163_ (.A1(\rvsingle.dp.rf.rf[21][18] ),
    .A2(_01296_),
    .B1(_01309_),
    .Y(_02084_));
 sky130_fd_sc_hd__o21a_2 _07164_ (.A1(_01432_),
    .A2(\rvsingle.dp.rf.rf[22][18] ),
    .B1(_01728_),
    .X(_02085_));
 sky130_fd_sc_hd__o21ai_2 _07165_ (.A1(\rvsingle.dp.rf.rf[23][18] ),
    .A2(_01943_),
    .B1(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__o211ai_2 _07166_ (.A1(_02083_),
    .A2(_02084_),
    .B1(_01703_),
    .C1(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__o211ai_2 _07167_ (.A1(_01915_),
    .A2(_02082_),
    .B1(_02087_),
    .C1(_01218_),
    .Y(_02088_));
 sky130_fd_sc_hd__or2_2 _07168_ (.A(_01417_),
    .B(\rvsingle.dp.rf.rf[24][18] ),
    .X(_02089_));
 sky130_fd_sc_hd__o211ai_2 _07169_ (.A1(\rvsingle.dp.rf.rf[25][18] ),
    .A2(_01943_),
    .B1(_01717_),
    .C1(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__o21a_2 _07170_ (.A1(_01242_),
    .A2(\rvsingle.dp.rf.rf[26][18] ),
    .B1(_01471_),
    .X(_02091_));
 sky130_fd_sc_hd__o21ai_2 _07171_ (.A1(\rvsingle.dp.rf.rf[27][18] ),
    .A2(_01943_),
    .B1(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__buf_1 _07172_ (.A(_01460_),
    .X(_02093_));
 sky130_fd_sc_hd__mux4_2 _07173_ (.A0(\rvsingle.dp.rf.rf[28][18] ),
    .A1(\rvsingle.dp.rf.rf[29][18] ),
    .A2(\rvsingle.dp.rf.rf[30][18] ),
    .A3(\rvsingle.dp.rf.rf[31][18] ),
    .S0(_01241_),
    .S1(_01199_),
    .X(_02094_));
 sky130_fd_sc_hd__o21ai_2 _07174_ (.A1(_02093_),
    .A2(_02094_),
    .B1(_01447_),
    .Y(_02095_));
 sky130_fd_sc_hd__a31o_2 _07175_ (.A1(_01208_),
    .A2(_02090_),
    .A3(_02092_),
    .B1(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__a31o_2 _07176_ (.A1(_02088_),
    .A2(_01450_),
    .A3(_02096_),
    .B1(_01452_),
    .X(_02097_));
 sky130_fd_sc_hd__o2bb2ai_2 _07177_ (.A1_N(_02066_),
    .A2_N(_02068_),
    .B1(_02081_),
    .B2(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__o211ai_2 _07178_ (.A1(_01223_),
    .A2(_02074_),
    .B1(_02080_),
    .C1(_01317_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand4b_2 _07179_ (.A_N(_02097_),
    .B(_02066_),
    .C(_02068_),
    .D(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__and4_2 _07180_ (.A(_02015_),
    .B(_02016_),
    .C(_02098_),
    .D(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__buf_1 _07181_ (.A(_01074_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_2 _07182_ (.A(_01666_),
    .B(\rvsingle.dp.rf.rf[26][17] ),
    .Y(_02103_));
 sky130_fd_sc_hd__o21ai_2 _07183_ (.A1(\rvsingle.dp.rf.rf[27][17] ),
    .A2(_01088_),
    .B1(_01626_),
    .Y(_02104_));
 sky130_fd_sc_hd__or2b_2 _07184_ (.A(\rvsingle.dp.rf.rf[25][17] ),
    .B_N(_01847_),
    .X(_02105_));
 sky130_fd_sc_hd__o211ai_2 _07185_ (.A1(_01848_),
    .A2(\rvsingle.dp.rf.rf[24][17] ),
    .B1(_02105_),
    .C1(_01759_),
    .Y(_02106_));
 sky130_fd_sc_hd__o21ai_2 _07186_ (.A1(_02103_),
    .A2(_02104_),
    .B1(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__nor2_2 _07187_ (.A(_01666_),
    .B(\rvsingle.dp.rf.rf[28][17] ),
    .Y(_02108_));
 sky130_fd_sc_hd__o21ai_2 _07188_ (.A1(\rvsingle.dp.rf.rf[29][17] ),
    .A2(_01842_),
    .B1(_01668_),
    .Y(_02109_));
 sky130_fd_sc_hd__o21a_2 _07189_ (.A1(_01763_),
    .A2(\rvsingle.dp.rf.rf[30][17] ),
    .B1(_01777_),
    .X(_02110_));
 sky130_fd_sc_hd__o21ai_2 _07190_ (.A1(\rvsingle.dp.rf.rf[31][17] ),
    .A2(_01861_),
    .B1(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__o211ai_2 _07191_ (.A1(_02108_),
    .A2(_02109_),
    .B1(_01503_),
    .C1(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__o211ai_2 _07192_ (.A1(_01512_),
    .A2(_02107_),
    .B1(_02112_),
    .C1(_01526_),
    .Y(_02113_));
 sky130_fd_sc_hd__o21bai_2 _07193_ (.A1(_01603_),
    .A2(\rvsingle.dp.rf.rf[16][17] ),
    .B1_N(_02031_),
    .Y(_02114_));
 sky130_fd_sc_hd__and2b_2 _07194_ (.A_N(\rvsingle.dp.rf.rf[17][17] ),
    .B(_01499_),
    .X(_02115_));
 sky130_fd_sc_hd__o21ai_2 _07195_ (.A1(_02114_),
    .A2(_02115_),
    .B1(_01565_),
    .Y(_02116_));
 sky130_fd_sc_hd__buf_1 _07196_ (.A(_01752_),
    .X(_02117_));
 sky130_fd_sc_hd__or2_2 _07197_ (.A(_02117_),
    .B(\rvsingle.dp.rf.rf[18][17] ),
    .X(_02118_));
 sky130_fd_sc_hd__o211a_2 _07198_ (.A1(_01865_),
    .A2(\rvsingle.dp.rf.rf[19][17] ),
    .B1(_01626_),
    .C1(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__nor2_2 _07199_ (.A(_01848_),
    .B(\rvsingle.dp.rf.rf[20][17] ),
    .Y(_02120_));
 sky130_fd_sc_hd__o21ai_2 _07200_ (.A1(\rvsingle.dp.rf.rf[21][17] ),
    .A2(_01842_),
    .B1(_01668_),
    .Y(_02121_));
 sky130_fd_sc_hd__o21a_2 _07201_ (.A1(_01763_),
    .A2(\rvsingle.dp.rf.rf[22][17] ),
    .B1(_01777_),
    .X(_02122_));
 sky130_fd_sc_hd__o21ai_2 _07202_ (.A1(\rvsingle.dp.rf.rf[23][17] ),
    .A2(_01861_),
    .B1(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__o211ai_2 _07203_ (.A1(_02120_),
    .A2(_02121_),
    .B1(_01503_),
    .C1(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__o211ai_2 _07204_ (.A1(_02116_),
    .A2(_02119_),
    .B1(_01634_),
    .C1(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__nand3_2 _07205_ (.A(_02113_),
    .B(_02125_),
    .C(_01682_),
    .Y(_02126_));
 sky130_fd_sc_hd__or2_2 _07206_ (.A(_01148_),
    .B(\rvsingle.dp.rf.rf[8][17] ),
    .X(_02127_));
 sky130_fd_sc_hd__o211a_2 _07207_ (.A1(\rvsingle.dp.rf.rf[9][17] ),
    .A2(_01088_),
    .B1(_01668_),
    .C1(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__nor2_2 _07208_ (.A(_01126_),
    .B(\rvsingle.dp.rf.rf[10][17] ),
    .Y(_02129_));
 sky130_fd_sc_hd__and2b_2 _07209_ (.A_N(\rvsingle.dp.rf.rf[11][17] ),
    .B(_02030_),
    .X(_02130_));
 sky130_fd_sc_hd__o31ai_2 _07210_ (.A1(_01759_),
    .A2(_02129_),
    .A3(_02130_),
    .B1(_01768_),
    .Y(_02131_));
 sky130_fd_sc_hd__o21ai_2 _07211_ (.A1(_01744_),
    .A2(\rvsingle.dp.rf.rf[14][17] ),
    .B1(_01648_),
    .Y(_02132_));
 sky130_fd_sc_hd__nor2_2 _07212_ (.A(\rvsingle.dp.rf.rf[15][17] ),
    .B(_01861_),
    .Y(_02133_));
 sky130_fd_sc_hd__or2_2 _07213_ (.A(_01753_),
    .B(\rvsingle.dp.rf.rf[12][17] ),
    .X(_02134_));
 sky130_fd_sc_hd__o211ai_2 _07214_ (.A1(\rvsingle.dp.rf.rf[13][17] ),
    .A2(_01865_),
    .B1(_01668_),
    .C1(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hd__o211ai_2 _07215_ (.A1(_02132_),
    .A2(_02133_),
    .B1(_01503_),
    .C1(_02135_),
    .Y(_02136_));
 sky130_fd_sc_hd__o211ai_2 _07216_ (.A1(_02128_),
    .A2(_02131_),
    .B1(_01526_),
    .C1(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_2 _07217_ (.A(_01666_),
    .B(\rvsingle.dp.rf.rf[6][17] ),
    .Y(_02138_));
 sky130_fd_sc_hd__o21ai_2 _07218_ (.A1(\rvsingle.dp.rf.rf[7][17] ),
    .A2(_01088_),
    .B1(_01626_),
    .Y(_02139_));
 sky130_fd_sc_hd__or2_2 _07219_ (.A(_01753_),
    .B(\rvsingle.dp.rf.rf[4][17] ),
    .X(_02140_));
 sky130_fd_sc_hd__o211ai_2 _07220_ (.A1(\rvsingle.dp.rf.rf[5][17] ),
    .A2(_01865_),
    .B1(_01668_),
    .C1(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__o211ai_2 _07221_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_01503_),
    .C1(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_2 _07222_ (.A(_01666_),
    .B(\rvsingle.dp.rf.rf[2][17] ),
    .Y(_02143_));
 sky130_fd_sc_hd__o21ai_2 _07223_ (.A1(\rvsingle.dp.rf.rf[3][17] ),
    .A2(_01088_),
    .B1(_01626_),
    .Y(_02144_));
 sky130_fd_sc_hd__or2_2 _07224_ (.A(_01607_),
    .B(\rvsingle.dp.rf.rf[0][17] ),
    .X(_02145_));
 sky130_fd_sc_hd__o211ai_2 _07225_ (.A1(\rvsingle.dp.rf.rf[1][17] ),
    .A2(_01842_),
    .B1(_01092_),
    .C1(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__o211ai_2 _07226_ (.A1(_02143_),
    .A2(_02144_),
    .B1(_02146_),
    .C1(_01565_),
    .Y(_02147_));
 sky130_fd_sc_hd__nand3_2 _07227_ (.A(_01634_),
    .B(_02142_),
    .C(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__nand3_2 _07228_ (.A(_01593_),
    .B(_02137_),
    .C(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__o211ai_2 _07229_ (.A1(_01962_),
    .A2(_01100_),
    .B1(_02126_),
    .C1(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__o221ai_2 _07230_ (.A1(_01960_),
    .A2(_02102_),
    .B1(_01961_),
    .B2(_02150_),
    .C1(_01587_),
    .Y(_02151_));
 sky130_fd_sc_hd__a31o_2 _07231_ (.A1(_01592_),
    .A2(_02149_),
    .A3(_02126_),
    .B1(_01178_),
    .X(_02152_));
 sky130_fd_sc_hd__o211ai_2 _07232_ (.A1(_01482_),
    .A2(_01171_),
    .B1(_01584_),
    .C1(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__mux4_2 _07233_ (.A0(\rvsingle.dp.rf.rf[0][17] ),
    .A1(\rvsingle.dp.rf.rf[1][17] ),
    .A2(\rvsingle.dp.rf.rf[2][17] ),
    .A3(\rvsingle.dp.rf.rf[3][17] ),
    .S0(_01726_),
    .S1(_01728_),
    .X(_02154_));
 sky130_fd_sc_hd__nor2_2 _07234_ (.A(_01703_),
    .B(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__mux2_2 _07235_ (.A0(\rvsingle.dp.rf.rf[4][17] ),
    .A1(\rvsingle.dp.rf.rf[5][17] ),
    .S(_01417_),
    .X(_02156_));
 sky130_fd_sc_hd__or2_2 _07236_ (.A(_01691_),
    .B(\rvsingle.dp.rf.rf[6][17] ),
    .X(_02157_));
 sky130_fd_sc_hd__o211a_2 _07237_ (.A1(_01688_),
    .A2(\rvsingle.dp.rf.rf[7][17] ),
    .B1(_01456_),
    .C1(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__a211oi_2 _07238_ (.A1(_02156_),
    .A2(_01717_),
    .B1(_01461_),
    .C1(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__mux4_2 _07239_ (.A0(\rvsingle.dp.rf.rf[12][17] ),
    .A1(\rvsingle.dp.rf.rf[13][17] ),
    .A2(\rvsingle.dp.rf.rf[14][17] ),
    .A3(\rvsingle.dp.rf.rf[15][17] ),
    .S0(_01192_),
    .S1(_01728_),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_2 _07240_ (.A0(\rvsingle.dp.rf.rf[8][17] ),
    .A1(\rvsingle.dp.rf.rf[9][17] ),
    .S(_01241_),
    .X(_02161_));
 sky130_fd_sc_hd__buf_1 _07241_ (.A(_01299_),
    .X(_02162_));
 sky130_fd_sc_hd__buf_1 _07242_ (.A(_01190_),
    .X(_02163_));
 sky130_fd_sc_hd__or2_2 _07243_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[10][17] ),
    .X(_02164_));
 sky130_fd_sc_hd__o211a_2 _07244_ (.A1(_01440_),
    .A2(\rvsingle.dp.rf.rf[11][17] ),
    .B1(_02162_),
    .C1(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__a211o_2 _07245_ (.A1(_02161_),
    .A2(_01437_),
    .B1(_01702_),
    .C1(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__o211ai_2 _07246_ (.A1(_01722_),
    .A2(_02160_),
    .B1(_01478_),
    .C1(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__o31ai_2 _07247_ (.A1(_01478_),
    .A2(_02155_),
    .A3(_02159_),
    .B1(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__mux2_2 _07248_ (.A0(\rvsingle.dp.rf.rf[28][17] ),
    .A1(\rvsingle.dp.rf.rf[29][17] ),
    .S(_01432_),
    .X(_02169_));
 sky130_fd_sc_hd__or2_2 _07249_ (.A(_01420_),
    .B(\rvsingle.dp.rf.rf[30][17] ),
    .X(_02170_));
 sky130_fd_sc_hd__o211a_2 _07250_ (.A1(_01688_),
    .A2(\rvsingle.dp.rf.rf[31][17] ),
    .B1(_01301_),
    .C1(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__a211oi_2 _07251_ (.A1(_02169_),
    .A2(_01717_),
    .B1(_01722_),
    .C1(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__mux4_2 _07252_ (.A0(\rvsingle.dp.rf.rf[24][17] ),
    .A1(\rvsingle.dp.rf.rf[25][17] ),
    .A2(\rvsingle.dp.rf.rf[26][17] ),
    .A3(\rvsingle.dp.rf.rf[27][17] ),
    .S0(_01469_),
    .S1(_01728_),
    .X(_02173_));
 sky130_fd_sc_hd__o21ai_2 _07253_ (.A1(_01703_),
    .A2(_02173_),
    .B1(_01478_),
    .Y(_02174_));
 sky130_fd_sc_hd__mux4_2 _07254_ (.A0(\rvsingle.dp.rf.rf[16][17] ),
    .A1(\rvsingle.dp.rf.rf[17][17] ),
    .A2(\rvsingle.dp.rf.rf[18][17] ),
    .A3(\rvsingle.dp.rf.rf[19][17] ),
    .S0(_01329_),
    .S1(_01456_),
    .X(_02175_));
 sky130_fd_sc_hd__buf_1 _07255_ (.A(_01425_),
    .X(_02176_));
 sky130_fd_sc_hd__mux4_2 _07256_ (.A0(\rvsingle.dp.rf.rf[20][17] ),
    .A1(\rvsingle.dp.rf.rf[21][17] ),
    .A2(\rvsingle.dp.rf.rf[22][17] ),
    .A3(\rvsingle.dp.rf.rf[23][17] ),
    .S0(_02176_),
    .S1(_01696_),
    .X(_02177_));
 sky130_fd_sc_hd__o21a_2 _07257_ (.A1(_02093_),
    .A2(_02177_),
    .B1(_01699_),
    .X(_02178_));
 sky130_fd_sc_hd__o21ai_2 _07258_ (.A1(_01230_),
    .A2(_02175_),
    .B1(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__o211ai_2 _07259_ (.A1(_02172_),
    .A2(_02174_),
    .B1(_01188_),
    .C1(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__o211a_2 _07260_ (.A1(_01450_),
    .A2(_02168_),
    .B1(_02180_),
    .C1(_01247_),
    .X(_02181_));
 sky130_fd_sc_hd__a21oi_2 _07261_ (.A1(_02151_),
    .A2(_02153_),
    .B1(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__nand3_2 _07262_ (.A(_02181_),
    .B(_02151_),
    .C(_02153_),
    .Y(_02183_));
 sky130_fd_sc_hd__nor2b_2 _07263_ (.A(_02182_),
    .B_N(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__o21a_2 _07264_ (.A1(_01336_),
    .A2(\rvsingle.dp.rf.rf[18][16] ),
    .B1(_01301_),
    .X(_02185_));
 sky130_fd_sc_hd__o21ai_2 _07265_ (.A1(\rvsingle.dp.rf.rf[19][16] ),
    .A2(_01943_),
    .B1(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__mux2_2 _07266_ (.A0(\rvsingle.dp.rf.rf[16][16] ),
    .A1(\rvsingle.dp.rf.rf[17][16] ),
    .S(_01417_),
    .X(_02187_));
 sky130_fd_sc_hd__a21oi_2 _07267_ (.A1(_02187_),
    .A2(_01717_),
    .B1(_01703_),
    .Y(_02188_));
 sky130_fd_sc_hd__mux4_2 _07268_ (.A0(\rvsingle.dp.rf.rf[20][16] ),
    .A1(\rvsingle.dp.rf.rf[21][16] ),
    .A2(\rvsingle.dp.rf.rf[22][16] ),
    .A3(\rvsingle.dp.rf.rf[23][16] ),
    .S0(_01432_),
    .S1(_01434_),
    .X(_02189_));
 sky130_fd_sc_hd__o2bb2ai_2 _07269_ (.A1_N(_02186_),
    .A2_N(_02188_),
    .B1(_01208_),
    .B2(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__buf_1 _07270_ (.A(_02093_),
    .X(_02191_));
 sky130_fd_sc_hd__mux4_2 _07271_ (.A0(\rvsingle.dp.rf.rf[28][16] ),
    .A1(\rvsingle.dp.rf.rf[29][16] ),
    .A2(\rvsingle.dp.rf.rf[30][16] ),
    .A3(\rvsingle.dp.rf.rf[31][16] ),
    .S0(_01242_),
    .S1(_01434_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_2 _07272_ (.A0(\rvsingle.dp.rf.rf[26][16] ),
    .A1(\rvsingle.dp.rf.rf[27][16] ),
    .S(_01726_),
    .X(_02193_));
 sky130_fd_sc_hd__or2_2 _07273_ (.A(_02176_),
    .B(\rvsingle.dp.rf.rf[24][16] ),
    .X(_02194_));
 sky130_fd_sc_hd__o211a_2 _07274_ (.A1(\rvsingle.dp.rf.rf[25][16] ),
    .A2(_01424_),
    .B1(_01716_),
    .C1(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__a211o_2 _07275_ (.A1(_01451_),
    .A2(_02193_),
    .B1(_02195_),
    .C1(_01445_),
    .X(_02196_));
 sky130_fd_sc_hd__o211ai_2 _07276_ (.A1(_02191_),
    .A2(_02192_),
    .B1(_01222_),
    .C1(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__o21ai_2 _07277_ (.A1(_01222_),
    .A2(_02190_),
    .B1(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__mux4_2 _07278_ (.A0(\rvsingle.dp.rf.rf[4][16] ),
    .A1(\rvsingle.dp.rf.rf[5][16] ),
    .A2(\rvsingle.dp.rf.rf[6][16] ),
    .A3(\rvsingle.dp.rf.rf[7][16] ),
    .S0(_01242_),
    .S1(_01200_),
    .X(_02199_));
 sky130_fd_sc_hd__or2_2 _07279_ (.A(_01469_),
    .B(\rvsingle.dp.rf.rf[0][16] ),
    .X(_02200_));
 sky130_fd_sc_hd__o211ai_2 _07280_ (.A1(\rvsingle.dp.rf.rf[1][16] ),
    .A2(_01296_),
    .B1(_01309_),
    .C1(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__o21a_2 _07281_ (.A1(_01417_),
    .A2(\rvsingle.dp.rf.rf[2][16] ),
    .B1(_01244_),
    .X(_02202_));
 sky130_fd_sc_hd__o21ai_2 _07282_ (.A1(\rvsingle.dp.rf.rf[3][16] ),
    .A2(_01296_),
    .B1(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__a31oi_2 _07283_ (.A1(_01722_),
    .A2(_02201_),
    .A3(_02203_),
    .B1(_01478_),
    .Y(_02204_));
 sky130_fd_sc_hd__o21ai_2 _07284_ (.A1(_02191_),
    .A2(_02199_),
    .B1(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__mux4_2 _07285_ (.A0(\rvsingle.dp.rf.rf[12][16] ),
    .A1(\rvsingle.dp.rf.rf[13][16] ),
    .A2(\rvsingle.dp.rf.rf[14][16] ),
    .A3(\rvsingle.dp.rf.rf[15][16] ),
    .S0(_01336_),
    .S1(_01200_),
    .X(_02206_));
 sky130_fd_sc_hd__mux4_2 _07286_ (.A0(\rvsingle.dp.rf.rf[8][16] ),
    .A1(\rvsingle.dp.rf.rf[9][16] ),
    .A2(\rvsingle.dp.rf.rf[10][16] ),
    .A3(\rvsingle.dp.rf.rf[11][16] ),
    .S0(_01707_),
    .S1(_01244_),
    .X(_02207_));
 sky130_fd_sc_hd__o21a_2 _07287_ (.A1(_01445_),
    .A2(_02207_),
    .B1(_01447_),
    .X(_02208_));
 sky130_fd_sc_hd__o21ai_2 _07288_ (.A1(_02191_),
    .A2(_02206_),
    .B1(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand3_2 _07289_ (.A(_01317_),
    .B(_02205_),
    .C(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__o211ai_2 _07290_ (.A1(_01317_),
    .A2(_02198_),
    .B1(_02210_),
    .C1(_01248_),
    .Y(_02211_));
 sky130_fd_sc_hd__clkdlybuf4s15_2 _07291_ (.A(_01128_),
    .X(_02212_));
 sky130_fd_sc_hd__nor2_2 _07292_ (.A(_01138_),
    .B(\rvsingle.dp.rf.rf[18][16] ),
    .Y(_02213_));
 sky130_fd_sc_hd__o21ai_2 _07293_ (.A1(\rvsingle.dp.rf.rf[19][16] ),
    .A2(_01509_),
    .B1(_01491_),
    .Y(_02214_));
 sky130_fd_sc_hd__or2_2 _07294_ (.A(_01595_),
    .B(\rvsingle.dp.rf.rf[16][16] ),
    .X(_02215_));
 sky130_fd_sc_hd__o211ai_2 _07295_ (.A1(\rvsingle.dp.rf.rf[17][16] ),
    .A2(_01488_),
    .B1(_01497_),
    .C1(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__o211a_2 _07296_ (.A1(_02213_),
    .A2(_02214_),
    .B1(_01132_),
    .C1(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__or2b_2 _07297_ (.A(\rvsingle.dp.rf.rf[21][16] ),
    .B_N(_01513_),
    .X(_02218_));
 sky130_fd_sc_hd__o211ai_2 _07298_ (.A1(_01269_),
    .A2(\rvsingle.dp.rf.rf[20][16] ),
    .B1(_02218_),
    .C1(_01497_),
    .Y(_02219_));
 sky130_fd_sc_hd__or2b_2 _07299_ (.A(\rvsingle.dp.rf.rf[23][16] ),
    .B_N(_01513_),
    .X(_02220_));
 sky130_fd_sc_hd__o211ai_2 _07300_ (.A1(_01383_),
    .A2(\rvsingle.dp.rf.rf[22][16] ),
    .B1(_01260_),
    .C1(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__a31o_2 _07301_ (.A1(_02219_),
    .A2(_02221_),
    .A3(_01512_),
    .B1(_01116_),
    .X(_02222_));
 sky130_fd_sc_hd__inv_2 _07302_ (.A(\rvsingle.dp.rf.rf[27][16] ),
    .Y(_02223_));
 sky130_fd_sc_hd__o21ai_2 _07303_ (.A1(_01098_),
    .A2(\rvsingle.dp.rf.rf[26][16] ),
    .B1(_01260_),
    .Y(_02224_));
 sky130_fd_sc_hd__a21oi_2 _07304_ (.A1(_02223_),
    .A2(_01257_),
    .B1(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__or2b_2 _07305_ (.A(\rvsingle.dp.rf.rf[25][16] ),
    .B_N(_02030_),
    .X(_02226_));
 sky130_fd_sc_hd__o211a_2 _07306_ (.A1(_01383_),
    .A2(\rvsingle.dp.rf.rf[24][16] ),
    .B1(_02226_),
    .C1(_01543_),
    .X(_02227_));
 sky130_fd_sc_hd__nor2_2 _07307_ (.A(_01383_),
    .B(\rvsingle.dp.rf.rf[28][16] ),
    .Y(_02228_));
 sky130_fd_sc_hd__o21ai_2 _07308_ (.A1(\rvsingle.dp.rf.rf[29][16] ),
    .A2(_01540_),
    .B1(_01543_),
    .Y(_02229_));
 sky130_fd_sc_hd__o21a_2 _07309_ (.A1(_01493_),
    .A2(\rvsingle.dp.rf.rf[30][16] ),
    .B1(_01523_),
    .X(_02230_));
 sky130_fd_sc_hd__o21ai_2 _07310_ (.A1(\rvsingle.dp.rf.rf[31][16] ),
    .A2(_01509_),
    .B1(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__o211ai_2 _07311_ (.A1(_02228_),
    .A2(_02229_),
    .B1(_01112_),
    .C1(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__o311ai_2 _07312_ (.A1(_01512_),
    .A2(_02225_),
    .A3(_02227_),
    .B1(_01506_),
    .C1(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__o211ai_2 _07313_ (.A1(_02217_),
    .A2(_02222_),
    .B1(_01147_),
    .C1(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__mux2_2 _07314_ (.A0(\rvsingle.dp.rf.rf[4][16] ),
    .A1(\rvsingle.dp.rf.rf[5][16] ),
    .S(_01666_),
    .X(_02235_));
 sky130_fd_sc_hd__buf_1 _07315_ (.A(_01768_),
    .X(_02236_));
 sky130_fd_sc_hd__or2b_2 _07316_ (.A(\rvsingle.dp.rf.rf[7][16] ),
    .B_N(_01518_),
    .X(_02237_));
 sky130_fd_sc_hd__o211a_2 _07317_ (.A1(_01269_),
    .A2(\rvsingle.dp.rf.rf[6][16] ),
    .B1(_01491_),
    .C1(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__a211oi_2 _07318_ (.A1(_02235_),
    .A2(_01093_),
    .B1(_02236_),
    .C1(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__or2_2 _07319_ (.A(_01595_),
    .B(\rvsingle.dp.rf.rf[2][16] ),
    .X(_02240_));
 sky130_fd_sc_hd__o211ai_2 _07320_ (.A1(_01488_),
    .A2(\rvsingle.dp.rf.rf[3][16] ),
    .B1(_01491_),
    .C1(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__or2b_2 _07321_ (.A(\rvsingle.dp.rf.rf[1][16] ),
    .B_N(_01595_),
    .X(_02242_));
 sky130_fd_sc_hd__o211ai_2 _07322_ (.A1(_01269_),
    .A2(\rvsingle.dp.rf.rf[0][16] ),
    .B1(_02242_),
    .C1(_01497_),
    .Y(_02243_));
 sky130_fd_sc_hd__a31o_2 _07323_ (.A1(_01132_),
    .A2(_02241_),
    .A3(_02243_),
    .B1(_01526_),
    .X(_02244_));
 sky130_fd_sc_hd__nor2_2 _07324_ (.A(_01269_),
    .B(\rvsingle.dp.rf.rf[14][16] ),
    .Y(_02245_));
 sky130_fd_sc_hd__o21ai_2 _07325_ (.A1(\rvsingle.dp.rf.rf[15][16] ),
    .A2(_01509_),
    .B1(_01491_),
    .Y(_02246_));
 sky130_fd_sc_hd__or2_2 _07326_ (.A(_01499_),
    .B(\rvsingle.dp.rf.rf[12][16] ),
    .X(_02247_));
 sky130_fd_sc_hd__o211ai_2 _07327_ (.A1(\rvsingle.dp.rf.rf[13][16] ),
    .A2(_01488_),
    .B1(_01543_),
    .C1(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__o21ai_2 _07328_ (.A1(_02245_),
    .A2(_02246_),
    .B1(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__nor2_2 _07329_ (.A(_01269_),
    .B(\rvsingle.dp.rf.rf[8][16] ),
    .Y(_02250_));
 sky130_fd_sc_hd__o21ai_2 _07330_ (.A1(\rvsingle.dp.rf.rf[9][16] ),
    .A2(_01509_),
    .B1(_01543_),
    .Y(_02251_));
 sky130_fd_sc_hd__o21a_2 _07331_ (.A1(_01562_),
    .A2(\rvsingle.dp.rf.rf[10][16] ),
    .B1(_01620_),
    .X(_02252_));
 sky130_fd_sc_hd__o21ai_2 _07332_ (.A1(\rvsingle.dp.rf.rf[11][16] ),
    .A2(_01488_),
    .B1(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__o211ai_2 _07333_ (.A1(_02250_),
    .A2(_02251_),
    .B1(_01132_),
    .C1(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__o211ai_2 _07334_ (.A1(_02236_),
    .A2(_02249_),
    .B1(_02254_),
    .C1(_01506_),
    .Y(_02255_));
 sky130_fd_sc_hd__o211ai_2 _07335_ (.A1(_02239_),
    .A2(_02244_),
    .B1(_01378_),
    .C1(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__o211ai_2 _07336_ (.A1(_01962_),
    .A2(_02212_),
    .B1(_02234_),
    .C1(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__a21oi_2 _07337_ (.A1(_02257_),
    .A2(_01482_),
    .B1(_01837_),
    .Y(_02258_));
 sky130_fd_sc_hd__buf_1 _07338_ (.A(Instr[4]),
    .X(_02259_));
 sky130_fd_sc_hd__nor4_2 _07339_ (.A(_02259_),
    .B(_01173_),
    .C(_01174_),
    .D(_01169_),
    .Y(_02260_));
 sky130_fd_sc_hd__o21ai_2 _07340_ (.A1(_01483_),
    .A2(_02260_),
    .B1(_01177_),
    .Y(_02261_));
 sky130_fd_sc_hd__nand4_2 _07341_ (.A(_02256_),
    .B(_01084_),
    .C(_01153_),
    .D(_02234_),
    .Y(_02262_));
 sky130_fd_sc_hd__o211a_2 _07342_ (.A1(_01066_),
    .A2(_01075_),
    .B1(_01587_),
    .C1(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__a21o_2 _07343_ (.A1(_02258_),
    .A2(_02261_),
    .B1(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__xor2_2 _07344_ (.A(_02211_),
    .B(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__nand4_2 _07345_ (.A(_01931_),
    .B(_02101_),
    .C(_02184_),
    .D(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__nor2_2 _07346_ (.A(_01695_),
    .B(\rvsingle.dp.rf.rf[12][7] ),
    .Y(_02267_));
 sky130_fd_sc_hd__buf_1 _07347_ (.A(_01306_),
    .X(_02268_));
 sky130_fd_sc_hd__o21ai_2 _07348_ (.A1(\rvsingle.dp.rf.rf[13][7] ),
    .A2(_01687_),
    .B1(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__nor2_2 _07349_ (.A(_01695_),
    .B(\rvsingle.dp.rf.rf[14][7] ),
    .Y(_02270_));
 sky130_fd_sc_hd__buf_1 _07350_ (.A(_01293_),
    .X(_02271_));
 sky130_fd_sc_hd__o21ai_2 _07351_ (.A1(\rvsingle.dp.rf.rf[15][7] ),
    .A2(_02271_),
    .B1(_01300_),
    .Y(_02272_));
 sky130_fd_sc_hd__buf_1 _07352_ (.A(_01172_),
    .X(_02273_));
 sky130_fd_sc_hd__o221a_2 _07353_ (.A1(_02267_),
    .A2(_02269_),
    .B1(_02270_),
    .B2(_02272_),
    .C1(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__buf_1 _07354_ (.A(_01294_),
    .X(_02275_));
 sky130_fd_sc_hd__o21ba_2 _07355_ (.A1(_01725_),
    .A2(\rvsingle.dp.rf.rf[8][7] ),
    .B1_N(_01299_),
    .X(_02276_));
 sky130_fd_sc_hd__o21ai_2 _07356_ (.A1(_02275_),
    .A2(\rvsingle.dp.rf.rf[9][7] ),
    .B1(_02276_),
    .Y(_02277_));
 sky130_fd_sc_hd__or2b_2 _07357_ (.A(\rvsingle.dp.rf.rf[11][7] ),
    .B_N(_02163_),
    .X(_02278_));
 sky130_fd_sc_hd__o211ai_2 _07358_ (.A1(_01420_),
    .A2(\rvsingle.dp.rf.rf[10][7] ),
    .B1(_01300_),
    .C1(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__a31o_2 _07359_ (.A1(_01460_),
    .A2(_02277_),
    .A3(_02279_),
    .B1(_01216_),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_2 _07360_ (.A0(\rvsingle.dp.rf.rf[0][7] ),
    .A1(\rvsingle.dp.rf.rf[1][7] ),
    .S(_01241_),
    .X(_02281_));
 sky130_fd_sc_hd__or2b_2 _07361_ (.A(\rvsingle.dp.rf.rf[3][7] ),
    .B_N(_01828_),
    .X(_02282_));
 sky130_fd_sc_hd__o211a_2 _07362_ (.A1(_01695_),
    .A2(\rvsingle.dp.rf.rf[2][7] ),
    .B1(_02162_),
    .C1(_02282_),
    .X(_02283_));
 sky130_fd_sc_hd__a211oi_2 _07363_ (.A1(_02281_),
    .A2(_01689_),
    .B1(_01702_),
    .C1(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__buf_1 _07364_ (.A(_01307_),
    .X(_02285_));
 sky130_fd_sc_hd__or2_2 _07365_ (.A(_01725_),
    .B(\rvsingle.dp.rf.rf[4][7] ),
    .X(_02286_));
 sky130_fd_sc_hd__o211ai_2 _07366_ (.A1(\rvsingle.dp.rf.rf[5][7] ),
    .A2(_01901_),
    .B1(_02285_),
    .C1(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__buf_1 _07367_ (.A(_01294_),
    .X(_02288_));
 sky130_fd_sc_hd__or2_2 _07368_ (.A(_01828_),
    .B(\rvsingle.dp.rf.rf[6][7] ),
    .X(_02289_));
 sky130_fd_sc_hd__o211ai_2 _07369_ (.A1(_02288_),
    .A2(\rvsingle.dp.rf.rf[7][7] ),
    .B1(_01808_),
    .C1(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__buf_1 _07370_ (.A(_01172_),
    .X(_02291_));
 sky130_fd_sc_hd__a31o_2 _07371_ (.A1(_02287_),
    .A2(_02290_),
    .A3(_02291_),
    .B1(_01446_),
    .X(_02292_));
 sky130_fd_sc_hd__o22ai_2 _07372_ (.A1(_02274_),
    .A2(_02280_),
    .B1(_02284_),
    .B2(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__mux4_2 _07373_ (.A0(\rvsingle.dp.rf.rf[28][7] ),
    .A1(\rvsingle.dp.rf.rf[29][7] ),
    .A2(\rvsingle.dp.rf.rf[30][7] ),
    .A3(\rvsingle.dp.rf.rf[31][7] ),
    .S0(_01426_),
    .S1(_01433_),
    .X(_02294_));
 sky130_fd_sc_hd__o21ai_2 _07374_ (.A1(_01192_),
    .A2(\rvsingle.dp.rf.rf[26][7] ),
    .B1(_01199_),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_2 _07375_ (.A(\rvsingle.dp.rf.rf[27][7] ),
    .B(_01424_),
    .Y(_02296_));
 sky130_fd_sc_hd__inv_2 _07376_ (.A(\rvsingle.dp.rf.rf[25][7] ),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_2 _07377_ (.A(_01416_),
    .B(\rvsingle.dp.rf.rf[24][7] ),
    .Y(_02298_));
 sky130_fd_sc_hd__a211o_2 _07378_ (.A1(_02297_),
    .A2(_01691_),
    .B1(_01727_),
    .C1(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__o211ai_2 _07379_ (.A1(_02295_),
    .A2(_02296_),
    .B1(_01721_),
    .C1(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__o211ai_2 _07380_ (.A1(_02093_),
    .A2(_02294_),
    .B1(_02300_),
    .C1(_01221_),
    .Y(_02301_));
 sky130_fd_sc_hd__buf_1 _07381_ (.A(_01444_),
    .X(_02302_));
 sky130_fd_sc_hd__buf_1 _07382_ (.A(_01294_),
    .X(_02303_));
 sky130_fd_sc_hd__or2_2 _07383_ (.A(_01468_),
    .B(\rvsingle.dp.rf.rf[18][7] ),
    .X(_02304_));
 sky130_fd_sc_hd__o211a_2 _07384_ (.A1(_02303_),
    .A2(\rvsingle.dp.rf.rf[19][7] ),
    .B1(_01953_),
    .C1(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__or2_2 _07385_ (.A(_01462_),
    .B(\rvsingle.dp.rf.rf[16][7] ),
    .X(_02306_));
 sky130_fd_sc_hd__o211a_2 _07386_ (.A1(\rvsingle.dp.rf.rf[17][7] ),
    .A2(_02303_),
    .B1(_02285_),
    .C1(_02306_),
    .X(_02307_));
 sky130_fd_sc_hd__inv_2 _07387_ (.A(\rvsingle.dp.rf.rf[21][7] ),
    .Y(_02308_));
 sky130_fd_sc_hd__nor2_2 _07388_ (.A(_01468_),
    .B(\rvsingle.dp.rf.rf[20][7] ),
    .Y(_02309_));
 sky130_fd_sc_hd__a211o_2 _07389_ (.A1(_02308_),
    .A2(_01730_),
    .B1(_01427_),
    .C1(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__o21a_2 _07390_ (.A1(_01725_),
    .A2(\rvsingle.dp.rf.rf[22][7] ),
    .B1(_01198_),
    .X(_02311_));
 sky130_fd_sc_hd__o21ai_2 _07391_ (.A1(\rvsingle.dp.rf.rf[23][7] ),
    .A2(_01827_),
    .B1(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__a31oi_2 _07392_ (.A1(_02310_),
    .A2(_02312_),
    .A3(_02291_),
    .B1(_01446_),
    .Y(_02313_));
 sky130_fd_sc_hd__o31ai_2 _07393_ (.A1(_02302_),
    .A2(_02305_),
    .A3(_02307_),
    .B1(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__buf_1 _07394_ (.A(Instr[19]),
    .X(_02315_));
 sky130_fd_sc_hd__nand3_2 _07395_ (.A(_02301_),
    .B(_02314_),
    .C(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__o211a_2 _07396_ (.A1(_01188_),
    .A2(_02293_),
    .B1(_02316_),
    .C1(_01246_),
    .X(_02317_));
 sky130_fd_sc_hd__buf_1 _07397_ (.A(_01074_),
    .X(_02318_));
 sky130_fd_sc_hd__inv_2 _07398_ (.A(Instr[27]),
    .Y(_02319_));
 sky130_fd_sc_hd__buf_1 _07399_ (.A(_01551_),
    .X(_02320_));
 sky130_fd_sc_hd__nor2_2 _07400_ (.A(_01862_),
    .B(\rvsingle.dp.rf.rf[12][7] ),
    .Y(_02321_));
 sky130_fd_sc_hd__and2b_2 _07401_ (.A_N(\rvsingle.dp.rf.rf[13][7] ),
    .B(_01618_),
    .X(_02322_));
 sky130_fd_sc_hd__buf_1 _07402_ (.A(_01110_),
    .X(_02323_));
 sky130_fd_sc_hd__or2b_2 _07403_ (.A(\rvsingle.dp.rf.rf[15][7] ),
    .B_N(_01544_),
    .X(_02324_));
 sky130_fd_sc_hd__o211ai_2 _07404_ (.A1(_01630_),
    .A2(\rvsingle.dp.rf.rf[14][7] ),
    .B1(_01259_),
    .C1(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__o311ai_2 _07405_ (.A1(_02320_),
    .A2(_02321_),
    .A3(_02322_),
    .B1(_02323_),
    .C1(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__nor2_2 _07406_ (.A(_01148_),
    .B(\rvsingle.dp.rf.rf[8][7] ),
    .Y(_02327_));
 sky130_fd_sc_hd__and2b_2 _07407_ (.A_N(\rvsingle.dp.rf.rf[9][7] ),
    .B(_01136_),
    .X(_02328_));
 sky130_fd_sc_hd__buf_1 _07408_ (.A(_01130_),
    .X(_02329_));
 sky130_fd_sc_hd__or2b_2 _07409_ (.A(\rvsingle.dp.rf.rf[11][7] ),
    .B_N(_01557_),
    .X(_02330_));
 sky130_fd_sc_hd__o211ai_2 _07410_ (.A1(_02117_),
    .A2(\rvsingle.dp.rf.rf[10][7] ),
    .B1(_01654_),
    .C1(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__o311ai_2 _07411_ (.A1(_01523_),
    .A2(_02327_),
    .A3(_02328_),
    .B1(_02329_),
    .C1(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__nand3_2 _07412_ (.A(_02326_),
    .B(_02332_),
    .C(_01505_),
    .Y(_02333_));
 sky130_fd_sc_hd__o21bai_2 _07413_ (.A1(_01753_),
    .A2(\rvsingle.dp.rf.rf[0][7] ),
    .B1_N(_01551_),
    .Y(_02334_));
 sky130_fd_sc_hd__and2b_2 _07414_ (.A_N(\rvsingle.dp.rf.rf[1][7] ),
    .B(_01618_),
    .X(_02335_));
 sky130_fd_sc_hd__o21ai_2 _07415_ (.A1(_02334_),
    .A2(_02335_),
    .B1(_02329_),
    .Y(_02336_));
 sky130_fd_sc_hd__buf_1 _07416_ (.A(_01519_),
    .X(_02337_));
 sky130_fd_sc_hd__or2b_2 _07417_ (.A(\rvsingle.dp.rf.rf[3][7] ),
    .B_N(_01498_),
    .X(_02338_));
 sky130_fd_sc_hd__o211a_2 _07418_ (.A1(_01780_),
    .A2(\rvsingle.dp.rf.rf[2][7] ),
    .B1(_02337_),
    .C1(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__nor2_2 _07419_ (.A(_02117_),
    .B(\rvsingle.dp.rf.rf[4][7] ),
    .Y(_02340_));
 sky130_fd_sc_hd__and2b_2 _07420_ (.A_N(\rvsingle.dp.rf.rf[5][7] ),
    .B(_01136_),
    .X(_02341_));
 sky130_fd_sc_hd__or2b_2 _07421_ (.A(\rvsingle.dp.rf.rf[7][7] ),
    .B_N(_01557_),
    .X(_02342_));
 sky130_fd_sc_hd__o211ai_2 _07422_ (.A1(_01658_),
    .A2(\rvsingle.dp.rf.rf[6][7] ),
    .B1(_01654_),
    .C1(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__o311ai_2 _07423_ (.A1(_01552_),
    .A2(_02340_),
    .A3(_02341_),
    .B1(_01111_),
    .C1(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__o211ai_2 _07424_ (.A1(_02336_),
    .A2(_02339_),
    .B1(_01156_),
    .C1(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand3_2 _07425_ (.A(_01377_),
    .B(_02333_),
    .C(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_2 _07426_ (.A(_01567_),
    .B(\rvsingle.dp.rf.rf[24][7] ),
    .Y(_02347_));
 sky130_fd_sc_hd__a211oi_2 _07427_ (.A1(_02297_),
    .A2(_01656_),
    .B1(_01620_),
    .C1(_02347_),
    .Y(_02348_));
 sky130_fd_sc_hd__o21ai_2 _07428_ (.A1(_01658_),
    .A2(\rvsingle.dp.rf.rf[26][7] ),
    .B1(_01259_),
    .Y(_02349_));
 sky130_fd_sc_hd__and2b_2 _07429_ (.A_N(\rvsingle.dp.rf.rf[27][7] ),
    .B(_01602_),
    .X(_02350_));
 sky130_fd_sc_hd__buf_1 _07430_ (.A(_01599_),
    .X(_02351_));
 sky130_fd_sc_hd__o21ai_2 _07431_ (.A1(_02349_),
    .A2(_02350_),
    .B1(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__nor2_2 _07432_ (.A(_01862_),
    .B(\rvsingle.dp.rf.rf[28][7] ),
    .Y(_02353_));
 sky130_fd_sc_hd__and2b_2 _07433_ (.A_N(\rvsingle.dp.rf.rf[29][7] ),
    .B(_01618_),
    .X(_02354_));
 sky130_fd_sc_hd__or2b_2 _07434_ (.A(\rvsingle.dp.rf.rf[31][7] ),
    .B_N(_01566_),
    .X(_02355_));
 sky130_fd_sc_hd__o211ai_2 _07435_ (.A1(_01630_),
    .A2(\rvsingle.dp.rf.rf[30][7] ),
    .B1(_01259_),
    .C1(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__o311ai_2 _07436_ (.A1(_02320_),
    .A2(_02353_),
    .A3(_02354_),
    .B1(_02323_),
    .C1(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__o211ai_2 _07437_ (.A1(_02348_),
    .A2(_02352_),
    .B1(_01505_),
    .C1(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__nor2_2 _07438_ (.A(_01630_),
    .B(\rvsingle.dp.rf.rf[20][7] ),
    .Y(_02359_));
 sky130_fd_sc_hd__a211oi_2 _07439_ (.A1(_02308_),
    .A2(_01614_),
    .B1(_02320_),
    .C1(_02359_),
    .Y(_02360_));
 sky130_fd_sc_hd__o21ai_2 _07440_ (.A1(_01675_),
    .A2(\rvsingle.dp.rf.rf[22][7] ),
    .B1(_01654_),
    .Y(_02361_));
 sky130_fd_sc_hd__and2b_2 _07441_ (.A_N(\rvsingle.dp.rf.rf[23][7] ),
    .B(_01561_),
    .X(_02362_));
 sky130_fd_sc_hd__o21ai_2 _07442_ (.A1(_02361_),
    .A2(_02362_),
    .B1(_02323_),
    .Y(_02363_));
 sky130_fd_sc_hd__buf_1 _07443_ (.A(_01155_),
    .X(_02364_));
 sky130_fd_sc_hd__nor2_2 _07444_ (.A(_02117_),
    .B(\rvsingle.dp.rf.rf[16][7] ),
    .Y(_02365_));
 sky130_fd_sc_hd__and2b_2 _07445_ (.A_N(\rvsingle.dp.rf.rf[17][7] ),
    .B(_01136_),
    .X(_02366_));
 sky130_fd_sc_hd__or2b_2 _07446_ (.A(\rvsingle.dp.rf.rf[19][7] ),
    .B_N(_01557_),
    .X(_02367_));
 sky130_fd_sc_hd__o211ai_2 _07447_ (.A1(_02117_),
    .A2(\rvsingle.dp.rf.rf[18][7] ),
    .B1(_01654_),
    .C1(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__o311ai_2 _07448_ (.A1(_01552_),
    .A2(_02365_),
    .A3(_02366_),
    .B1(_02329_),
    .C1(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__o211ai_2 _07449_ (.A1(_02360_),
    .A2(_02363_),
    .B1(_02364_),
    .C1(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__nand3_2 _07450_ (.A(_02358_),
    .B(_02370_),
    .C(_01146_),
    .Y(_02371_));
 sky130_fd_sc_hd__nand4_2 _07451_ (.A(_01152_),
    .B(_02346_),
    .C(_02371_),
    .D(_01083_),
    .Y(_02372_));
 sky130_fd_sc_hd__o221ai_2 _07452_ (.A1(_01065_),
    .A2(_02318_),
    .B1(_01870_),
    .B2(_02319_),
    .C1(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_2 _07453_ (.A(_02317_),
    .B(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__buf_1 _07454_ (.A(_01177_),
    .X(_02375_));
 sky130_fd_sc_hd__nand2_2 _07455_ (.A(_02375_),
    .B(Instr[27]),
    .Y(_02376_));
 sky130_fd_sc_hd__a21oi_2 _07456_ (.A1(_02376_),
    .A2(_02372_),
    .B1(_01485_),
    .Y(_02377_));
 sky130_fd_sc_hd__nor2_2 _07457_ (.A(_01763_),
    .B(\rvsingle.dp.rf.rf[26][6] ),
    .Y(_02378_));
 sky130_fd_sc_hd__buf_1 _07458_ (.A(_01086_),
    .X(_02379_));
 sky130_fd_sc_hd__o21ai_2 _07459_ (.A1(\rvsingle.dp.rf.rf[27][6] ),
    .A2(_02379_),
    .B1(_01777_),
    .Y(_02380_));
 sky130_fd_sc_hd__nor2_2 _07460_ (.A(_02030_),
    .B(\rvsingle.dp.rf.rf[24][6] ),
    .Y(_02381_));
 sky130_fd_sc_hd__o21ai_2 _07461_ (.A1(\rvsingle.dp.rf.rf[25][6] ),
    .A2(_01539_),
    .B1(_01542_),
    .Y(_02382_));
 sky130_fd_sc_hd__o221ai_2 _07462_ (.A1(_02378_),
    .A2(_02380_),
    .B1(_02381_),
    .B2(_02382_),
    .C1(_02351_),
    .Y(_02383_));
 sky130_fd_sc_hd__nor2_2 _07463_ (.A(_02117_),
    .B(\rvsingle.dp.rf.rf[30][6] ),
    .Y(_02384_));
 sky130_fd_sc_hd__and2b_2 _07464_ (.A_N(\rvsingle.dp.rf.rf[31][6] ),
    .B(_01613_),
    .X(_02385_));
 sky130_fd_sc_hd__o21ba_2 _07465_ (.A1(_01779_),
    .A2(\rvsingle.dp.rf.rf[28][6] ),
    .B1_N(_01610_),
    .X(_02386_));
 sky130_fd_sc_hd__o21ai_2 _07466_ (.A1(_02379_),
    .A2(\rvsingle.dp.rf.rf[29][6] ),
    .B1(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__o311ai_2 _07467_ (.A1(_01496_),
    .A2(_02384_),
    .A3(_02385_),
    .B1(_02323_),
    .C1(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__nand3_2 _07468_ (.A(_02383_),
    .B(_01505_),
    .C(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__nor2_2 _07469_ (.A(_01847_),
    .B(\rvsingle.dp.rf.rf[16][6] ),
    .Y(_02390_));
 sky130_fd_sc_hd__and2b_2 _07470_ (.A_N(\rvsingle.dp.rf.rf[17][6] ),
    .B(_01594_),
    .X(_02391_));
 sky130_fd_sc_hd__or2b_2 _07471_ (.A(\rvsingle.dp.rf.rf[19][6] ),
    .B_N(_01096_),
    .X(_02392_));
 sky130_fd_sc_hd__o211ai_2 _07472_ (.A1(_01675_),
    .A2(\rvsingle.dp.rf.rf[18][6] ),
    .B1(_01611_),
    .C1(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__o311ai_2 _07473_ (.A1(_01490_),
    .A2(_02390_),
    .A3(_02391_),
    .B1(_01564_),
    .C1(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__buf_1 _07474_ (.A(_01091_),
    .X(_02395_));
 sky130_fd_sc_hd__nor2_2 _07475_ (.A(_01847_),
    .B(\rvsingle.dp.rf.rf[22][6] ),
    .Y(_02396_));
 sky130_fd_sc_hd__and2b_2 _07476_ (.A_N(\rvsingle.dp.rf.rf[23][6] ),
    .B(_01594_),
    .X(_02397_));
 sky130_fd_sc_hd__o21ba_2 _07477_ (.A1(_01544_),
    .A2(\rvsingle.dp.rf.rf[20][6] ),
    .B1_N(_01610_),
    .X(_02398_));
 sky130_fd_sc_hd__o21ai_2 _07478_ (.A1(_01860_),
    .A2(\rvsingle.dp.rf.rf[21][6] ),
    .B1(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__o311ai_2 _07479_ (.A1(_02395_),
    .A2(_02396_),
    .A3(_02397_),
    .B1(_01111_),
    .C1(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand3_2 _07480_ (.A(_01156_),
    .B(_02394_),
    .C(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand3_2 _07481_ (.A(_02389_),
    .B(_02401_),
    .C(_01146_),
    .Y(_02402_));
 sky130_fd_sc_hd__or2b_2 _07482_ (.A(\rvsingle.dp.rf.rf[11][6] ),
    .B_N(_01877_),
    .X(_02403_));
 sky130_fd_sc_hd__o211a_2 _07483_ (.A1(_01763_),
    .A2(\rvsingle.dp.rf.rf[10][6] ),
    .B1(_02031_),
    .C1(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__o21bai_2 _07484_ (.A1(_01847_),
    .A2(\rvsingle.dp.rf.rf[8][6] ),
    .B1_N(_01551_),
    .Y(_02405_));
 sky130_fd_sc_hd__and2b_2 _07485_ (.A_N(\rvsingle.dp.rf.rf[9][6] ),
    .B(_01561_),
    .X(_02406_));
 sky130_fd_sc_hd__o21ai_2 _07486_ (.A1(_02405_),
    .A2(_02406_),
    .B1(_01131_),
    .Y(_02407_));
 sky130_fd_sc_hd__nor2_2 _07487_ (.A(_01545_),
    .B(\rvsingle.dp.rf.rf[12][6] ),
    .Y(_02408_));
 sky130_fd_sc_hd__o21ai_2 _07488_ (.A1(\rvsingle.dp.rf.rf[13][6] ),
    .A2(_02379_),
    .B1(_01542_),
    .Y(_02409_));
 sky130_fd_sc_hd__buf_1 _07489_ (.A(_01110_),
    .X(_02410_));
 sky130_fd_sc_hd__o21a_2 _07490_ (.A1(_01267_),
    .A2(\rvsingle.dp.rf.rf[14][6] ),
    .B1(_01489_),
    .X(_02411_));
 sky130_fd_sc_hd__o21ai_2 _07491_ (.A1(\rvsingle.dp.rf.rf[15][6] ),
    .A2(_01508_),
    .B1(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__o211ai_2 _07492_ (.A1(_02408_),
    .A2(_02409_),
    .B1(_02410_),
    .C1(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__o211ai_2 _07493_ (.A1(_02404_),
    .A2(_02407_),
    .B1(_01505_),
    .C1(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__nor2_2 _07494_ (.A(_02117_),
    .B(\rvsingle.dp.rf.rf[0][6] ),
    .Y(_02415_));
 sky130_fd_sc_hd__and2b_2 _07495_ (.A_N(\rvsingle.dp.rf.rf[1][6] ),
    .B(_01613_),
    .X(_02416_));
 sky130_fd_sc_hd__or2b_2 _07496_ (.A(\rvsingle.dp.rf.rf[3][6] ),
    .B_N(_01557_),
    .X(_02417_));
 sky130_fd_sc_hd__o211ai_2 _07497_ (.A1(_01658_),
    .A2(\rvsingle.dp.rf.rf[2][6] ),
    .B1(_01654_),
    .C1(_02417_),
    .Y(_02418_));
 sky130_fd_sc_hd__o311ai_2 _07498_ (.A1(_01552_),
    .A2(_02415_),
    .A3(_02416_),
    .B1(_02329_),
    .C1(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__nor2_2 _07499_ (.A(_01097_),
    .B(\rvsingle.dp.rf.rf[4][6] ),
    .Y(_02420_));
 sky130_fd_sc_hd__and2b_2 _07500_ (.A_N(\rvsingle.dp.rf.rf[5][6] ),
    .B(_01613_),
    .X(_02421_));
 sky130_fd_sc_hd__or2b_2 _07501_ (.A(\rvsingle.dp.rf.rf[7][6] ),
    .B_N(_01557_),
    .X(_02422_));
 sky130_fd_sc_hd__o211ai_2 _07502_ (.A1(_01658_),
    .A2(\rvsingle.dp.rf.rf[6][6] ),
    .B1(_01654_),
    .C1(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__o311ai_2 _07503_ (.A1(_01552_),
    .A2(_02420_),
    .A3(_02421_),
    .B1(_02323_),
    .C1(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand3_2 _07504_ (.A(_01156_),
    .B(_02419_),
    .C(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__nand3_2 _07505_ (.A(_01377_),
    .B(_02414_),
    .C(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__o211ai_2 _07506_ (.A1(_01139_),
    .A2(_01962_),
    .B1(_02402_),
    .C1(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__nand2_2 _07507_ (.A(_02427_),
    .B(_01870_),
    .Y(_02428_));
 sky130_fd_sc_hd__or2_2 _07508_ (.A(Instr[26]),
    .B(_01083_),
    .X(_02429_));
 sky130_fd_sc_hd__nand3_2 _07509_ (.A(_02428_),
    .B(_01183_),
    .C(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__nand2_2 _07510_ (.A(_02375_),
    .B(Instr[26]),
    .Y(_02431_));
 sky130_fd_sc_hd__o221ai_2 _07511_ (.A1(_01065_),
    .A2(_02318_),
    .B1(_01178_),
    .B2(_02427_),
    .C1(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__mux2_2 _07512_ (.A0(\rvsingle.dp.rf.rf[8][6] ),
    .A1(\rvsingle.dp.rf.rf[9][6] ),
    .S(_01730_),
    .X(_02433_));
 sky130_fd_sc_hd__or2_2 _07513_ (.A(_01349_),
    .B(\rvsingle.dp.rf.rf[10][6] ),
    .X(_02434_));
 sky130_fd_sc_hd__o211a_2 _07514_ (.A1(_01440_),
    .A2(\rvsingle.dp.rf.rf[11][6] ),
    .B1(_01696_),
    .C1(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__a211oi_2 _07515_ (.A1(_02433_),
    .A2(_01689_),
    .B1(_01702_),
    .C1(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__mux4_2 _07516_ (.A0(\rvsingle.dp.rf.rf[12][6] ),
    .A1(\rvsingle.dp.rf.rf[13][6] ),
    .A2(\rvsingle.dp.rf.rf[14][6] ),
    .A3(\rvsingle.dp.rf.rf[15][6] ),
    .S0(_01462_),
    .S1(_01727_),
    .X(_02437_));
 sky130_fd_sc_hd__buf_1 _07517_ (.A(_01215_),
    .X(_02438_));
 sky130_fd_sc_hd__o21ai_2 _07518_ (.A1(_01207_),
    .A2(_02437_),
    .B1(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__buf_1 _07519_ (.A(_01327_),
    .X(_02440_));
 sky130_fd_sc_hd__mux4_2 _07520_ (.A0(\rvsingle.dp.rf.rf[0][6] ),
    .A1(\rvsingle.dp.rf.rf[1][6] ),
    .A2(\rvsingle.dp.rf.rf[2][6] ),
    .A3(\rvsingle.dp.rf.rf[3][6] ),
    .S0(_02440_),
    .S1(_01470_),
    .X(_02441_));
 sky130_fd_sc_hd__nor2_2 _07521_ (.A(_01707_),
    .B(\rvsingle.dp.rf.rf[4][6] ),
    .Y(_02442_));
 sky130_fd_sc_hd__o21ai_2 _07522_ (.A1(\rvsingle.dp.rf.rf[5][6] ),
    .A2(_01687_),
    .B1(_02268_),
    .Y(_02443_));
 sky130_fd_sc_hd__nor2_2 _07523_ (.A(_01707_),
    .B(\rvsingle.dp.rf.rf[6][6] ),
    .Y(_02444_));
 sky130_fd_sc_hd__o21ai_2 _07524_ (.A1(\rvsingle.dp.rf.rf[7][6] ),
    .A2(_01687_),
    .B1(_01708_),
    .Y(_02445_));
 sky130_fd_sc_hd__o221ai_2 _07525_ (.A1(_02442_),
    .A2(_02443_),
    .B1(_02444_),
    .B2(_02445_),
    .C1(_02273_),
    .Y(_02446_));
 sky130_fd_sc_hd__buf_1 _07526_ (.A(_01216_),
    .X(_02447_));
 sky130_fd_sc_hd__o211ai_2 _07527_ (.A1(_01229_),
    .A2(_02441_),
    .B1(_02446_),
    .C1(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__o21ai_2 _07528_ (.A1(_02436_),
    .A2(_02439_),
    .B1(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__buf_1 _07529_ (.A(_01327_),
    .X(_02450_));
 sky130_fd_sc_hd__mux4_2 _07530_ (.A0(\rvsingle.dp.rf.rf[24][6] ),
    .A1(\rvsingle.dp.rf.rf[25][6] ),
    .A2(\rvsingle.dp.rf.rf[26][6] ),
    .A3(\rvsingle.dp.rf.rf[27][6] ),
    .S0(_02450_),
    .S1(_01455_),
    .X(_02451_));
 sky130_fd_sc_hd__nor2_2 _07531_ (.A(_02302_),
    .B(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__mux4_2 _07532_ (.A0(\rvsingle.dp.rf.rf[28][6] ),
    .A1(\rvsingle.dp.rf.rf[29][6] ),
    .A2(\rvsingle.dp.rf.rf[30][6] ),
    .A3(\rvsingle.dp.rf.rf[31][6] ),
    .S0(_01462_),
    .S1(_01470_),
    .X(_02453_));
 sky130_fd_sc_hd__o21ai_2 _07533_ (.A1(_01207_),
    .A2(_02453_),
    .B1(_02438_),
    .Y(_02454_));
 sky130_fd_sc_hd__mux4_2 _07534_ (.A0(\rvsingle.dp.rf.rf[16][6] ),
    .A1(\rvsingle.dp.rf.rf[17][6] ),
    .A2(\rvsingle.dp.rf.rf[18][6] ),
    .A3(\rvsingle.dp.rf.rf[19][6] ),
    .S0(_01462_),
    .S1(_01727_),
    .X(_02455_));
 sky130_fd_sc_hd__nor2_2 _07535_ (.A(_01420_),
    .B(\rvsingle.dp.rf.rf[20][6] ),
    .Y(_02456_));
 sky130_fd_sc_hd__o21ai_2 _07536_ (.A1(\rvsingle.dp.rf.rf[21][6] ),
    .A2(_02271_),
    .B1(_02268_),
    .Y(_02457_));
 sky130_fd_sc_hd__o21a_2 _07537_ (.A1(_01725_),
    .A2(\rvsingle.dp.rf.rf[22][6] ),
    .B1(_01198_),
    .X(_02458_));
 sky130_fd_sc_hd__o21ai_2 _07538_ (.A1(\rvsingle.dp.rf.rf[23][6] ),
    .A2(_02288_),
    .B1(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__o211ai_2 _07539_ (.A1(_02456_),
    .A2(_02457_),
    .B1(_01444_),
    .C1(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__o211ai_2 _07540_ (.A1(_01229_),
    .A2(_02455_),
    .B1(_02460_),
    .C1(_02447_),
    .Y(_02461_));
 sky130_fd_sc_hd__o211ai_2 _07541_ (.A1(_02452_),
    .A2(_02454_),
    .B1(_02461_),
    .C1(_01187_),
    .Y(_02462_));
 sky130_fd_sc_hd__o211a_2 _07542_ (.A1(_02315_),
    .A2(_02449_),
    .B1(_02462_),
    .C1(_01246_),
    .X(_02463_));
 sky130_fd_sc_hd__nand3_2 _07543_ (.A(_02430_),
    .B(_02432_),
    .C(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__o21ai_2 _07544_ (.A1(_01450_),
    .A2(_02293_),
    .B1(_01247_),
    .Y(_02465_));
 sky130_fd_sc_hd__and3_2 _07545_ (.A(_02301_),
    .B(_02314_),
    .C(_01188_),
    .X(_02466_));
 sky130_fd_sc_hd__o221a_2 _07546_ (.A1(_01065_),
    .A2(_01074_),
    .B1(_01870_),
    .B2(_02319_),
    .C1(_02372_),
    .X(_02467_));
 sky130_fd_sc_hd__o22ai_2 _07547_ (.A1(_02465_),
    .A2(_02466_),
    .B1(_02467_),
    .B2(_02377_),
    .Y(_02468_));
 sky130_fd_sc_hd__buf_1 _07548_ (.A(_01452_),
    .X(_02469_));
 sky130_fd_sc_hd__o21ai_2 _07549_ (.A1(_01450_),
    .A2(_02449_),
    .B1(_02462_),
    .Y(_02470_));
 sky130_fd_sc_hd__nand4_2 _07550_ (.A(_01592_),
    .B(_02402_),
    .C(_02426_),
    .D(_01481_),
    .Y(_02471_));
 sky130_fd_sc_hd__a21oi_2 _07551_ (.A1(_02471_),
    .A2(_02431_),
    .B1(_01591_),
    .Y(_02472_));
 sky130_fd_sc_hd__buf_1 _07552_ (.A(_01064_),
    .X(_02473_));
 sky130_fd_sc_hd__o211a_2 _07553_ (.A1(_02473_),
    .A2(_02102_),
    .B1(_02471_),
    .C1(_02431_),
    .X(_02474_));
 sky130_fd_sc_hd__o22ai_2 _07554_ (.A1(_02469_),
    .A2(_02470_),
    .B1(_02472_),
    .B2(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__o2111a_2 _07555_ (.A1(_02374_),
    .A2(_02377_),
    .B1(_02464_),
    .C1(_02468_),
    .D1(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__nor2_2 _07556_ (.A(_01518_),
    .B(\rvsingle.dp.rf.rf[2][4] ),
    .Y(_02477_));
 sky130_fd_sc_hd__buf_1 _07557_ (.A(_01086_),
    .X(_02478_));
 sky130_fd_sc_hd__o21ai_2 _07558_ (.A1(\rvsingle.dp.rf.rf[3][4] ),
    .A2(_02478_),
    .B1(_01523_),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_2 _07559_ (.A(_01619_),
    .B(\rvsingle.dp.rf.rf[0][4] ),
    .Y(_02480_));
 sky130_fd_sc_hd__buf_1 _07560_ (.A(_01645_),
    .X(_02481_));
 sky130_fd_sc_hd__o21ai_2 _07561_ (.A1(\rvsingle.dp.rf.rf[1][4] ),
    .A2(_02481_),
    .B1(_01496_),
    .Y(_02482_));
 sky130_fd_sc_hd__buf_1 _07562_ (.A(_01599_),
    .X(_02483_));
 sky130_fd_sc_hd__o221a_2 _07563_ (.A1(_02477_),
    .A2(_02479_),
    .B1(_02480_),
    .B2(_02482_),
    .C1(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__buf_1 _07564_ (.A(_01091_),
    .X(_02485_));
 sky130_fd_sc_hd__or2_2 _07565_ (.A(_01136_),
    .B(\rvsingle.dp.rf.rf[4][4] ),
    .X(_02486_));
 sky130_fd_sc_hd__o211ai_2 _07566_ (.A1(\rvsingle.dp.rf.rf[5][4] ),
    .A2(_01677_),
    .B1(_02485_),
    .C1(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__buf_1 _07567_ (.A(_01110_),
    .X(_02488_));
 sky130_fd_sc_hd__or2b_2 _07568_ (.A(\rvsingle.dp.rf.rf[7][4] ),
    .B_N(_01618_),
    .X(_02489_));
 sky130_fd_sc_hd__o211ai_2 _07569_ (.A1(_01493_),
    .A2(\rvsingle.dp.rf.rf[6][4] ),
    .B1(_01552_),
    .C1(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__buf_1 _07570_ (.A(_01115_),
    .X(_02491_));
 sky130_fd_sc_hd__a31o_2 _07571_ (.A1(_02487_),
    .A2(_02488_),
    .A3(_02490_),
    .B1(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__nor2_2 _07572_ (.A(_01493_),
    .B(\rvsingle.dp.rf.rf[10][4] ),
    .Y(_02493_));
 sky130_fd_sc_hd__o21ai_2 _07573_ (.A1(\rvsingle.dp.rf.rf[11][4] ),
    .A2(_02478_),
    .B1(_01523_),
    .Y(_02494_));
 sky130_fd_sc_hd__o21ba_2 _07574_ (.A1(_01561_),
    .A2(\rvsingle.dp.rf.rf[8][4] ),
    .B1_N(_01489_),
    .X(_02495_));
 sky130_fd_sc_hd__o21ai_2 _07575_ (.A1(_02481_),
    .A2(\rvsingle.dp.rf.rf[9][4] ),
    .B1(_02495_),
    .Y(_02496_));
 sky130_fd_sc_hd__o21ai_2 _07576_ (.A1(_02493_),
    .A2(_02494_),
    .B1(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__nor2_2 _07577_ (.A(_01780_),
    .B(\rvsingle.dp.rf.rf[14][4] ),
    .Y(_02498_));
 sky130_fd_sc_hd__o21ai_2 _07578_ (.A1(\rvsingle.dp.rf.rf[15][4] ),
    .A2(_01539_),
    .B1(_01520_),
    .Y(_02499_));
 sky130_fd_sc_hd__nor2_2 _07579_ (.A(_01878_),
    .B(\rvsingle.dp.rf.rf[12][4] ),
    .Y(_02500_));
 sky130_fd_sc_hd__o21ai_2 _07580_ (.A1(\rvsingle.dp.rf.rf[13][4] ),
    .A2(_01508_),
    .B1(_02395_),
    .Y(_02501_));
 sky130_fd_sc_hd__o221ai_2 _07581_ (.A1(_02498_),
    .A2(_02499_),
    .B1(_02500_),
    .B2(_02501_),
    .C1(_02488_),
    .Y(_02502_));
 sky130_fd_sc_hd__o211ai_2 _07582_ (.A1(_01503_),
    .A2(_02497_),
    .B1(_02502_),
    .C1(_01116_),
    .Y(_02503_));
 sky130_fd_sc_hd__o211ai_2 _07583_ (.A1(_02484_),
    .A2(_02492_),
    .B1(_01377_),
    .C1(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__buf_1 _07584_ (.A(_01152_),
    .X(_02505_));
 sky130_fd_sc_hd__nor2_2 _07585_ (.A(_01518_),
    .B(\rvsingle.dp.rf.rf[18][4] ),
    .Y(_02506_));
 sky130_fd_sc_hd__o21ai_2 _07586_ (.A1(\rvsingle.dp.rf.rf[19][4] ),
    .A2(_02481_),
    .B1(_01552_),
    .Y(_02507_));
 sky130_fd_sc_hd__or2b_2 _07587_ (.A(\rvsingle.dp.rf.rf[17][4] ),
    .B_N(_01267_),
    .X(_02508_));
 sky130_fd_sc_hd__o211ai_2 _07588_ (.A1(_01513_),
    .A2(\rvsingle.dp.rf.rf[16][4] ),
    .B1(_02508_),
    .C1(_01496_),
    .Y(_02509_));
 sky130_fd_sc_hd__o211ai_2 _07589_ (.A1(_02506_),
    .A2(_02507_),
    .B1(_02509_),
    .C1(_01600_),
    .Y(_02510_));
 sky130_fd_sc_hd__nor2_2 _07590_ (.A(_01518_),
    .B(\rvsingle.dp.rf.rf[22][4] ),
    .Y(_02511_));
 sky130_fd_sc_hd__o21ai_2 _07591_ (.A1(\rvsingle.dp.rf.rf[23][4] ),
    .A2(_02481_),
    .B1(_02320_),
    .Y(_02512_));
 sky130_fd_sc_hd__or2b_2 _07592_ (.A(\rvsingle.dp.rf.rf[21][4] ),
    .B_N(_01267_),
    .X(_02513_));
 sky130_fd_sc_hd__o211ai_2 _07593_ (.A1(_01513_),
    .A2(\rvsingle.dp.rf.rf[20][4] ),
    .B1(_02513_),
    .C1(_02485_),
    .Y(_02514_));
 sky130_fd_sc_hd__o211ai_2 _07594_ (.A1(_02511_),
    .A2(_02512_),
    .B1(_02514_),
    .C1(_01617_),
    .Y(_02515_));
 sky130_fd_sc_hd__nand3_2 _07595_ (.A(_01853_),
    .B(_02510_),
    .C(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__nor2_2 _07596_ (.A(_01614_),
    .B(\rvsingle.dp.rf.rf[30][4] ),
    .Y(_02517_));
 sky130_fd_sc_hd__o21ai_2 _07597_ (.A1(\rvsingle.dp.rf.rf[31][4] ),
    .A2(_02481_),
    .B1(_02320_),
    .Y(_02518_));
 sky130_fd_sc_hd__or2b_2 _07598_ (.A(\rvsingle.dp.rf.rf[29][4] ),
    .B_N(_01267_),
    .X(_02519_));
 sky130_fd_sc_hd__o211ai_2 _07599_ (.A1(_01595_),
    .A2(\rvsingle.dp.rf.rf[28][4] ),
    .B1(_02519_),
    .C1(_02485_),
    .Y(_02520_));
 sky130_fd_sc_hd__o211ai_2 _07600_ (.A1(_02517_),
    .A2(_02518_),
    .B1(_02520_),
    .C1(_01617_),
    .Y(_02521_));
 sky130_fd_sc_hd__nor2_2 _07601_ (.A(_02030_),
    .B(\rvsingle.dp.rf.rf[24][4] ),
    .Y(_02522_));
 sky130_fd_sc_hd__and2b_2 _07602_ (.A_N(\rvsingle.dp.rf.rf[25][4] ),
    .B(_01602_),
    .X(_02523_));
 sky130_fd_sc_hd__o21a_2 _07603_ (.A1(_01136_),
    .A2(\rvsingle.dp.rf.rf[26][4] ),
    .B1(_01551_),
    .X(_02524_));
 sky130_fd_sc_hd__o21ai_2 _07604_ (.A1(\rvsingle.dp.rf.rf[27][4] ),
    .A2(_01487_),
    .B1(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__o311ai_2 _07605_ (.A1(_01660_),
    .A2(_02522_),
    .A3(_02523_),
    .B1(_02351_),
    .C1(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__buf_1 _07606_ (.A(_01115_),
    .X(_02527_));
 sky130_fd_sc_hd__nand3_2 _07607_ (.A(_02521_),
    .B(_02526_),
    .C(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__nand3_2 _07608_ (.A(_02516_),
    .B(_01146_),
    .C(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__nand4_2 _07609_ (.A(_02504_),
    .B(_01083_),
    .C(_02505_),
    .D(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__a31o_2 _07610_ (.A1(_01076_),
    .A2(_01071_),
    .A3(_01062_),
    .B1(_01145_),
    .X(_02531_));
 sky130_fd_sc_hd__o21a_2 _07611_ (.A1(Instr[11]),
    .A2(_01078_),
    .B1(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__nand2_2 _07612_ (.A(_01178_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__a21oi_2 _07613_ (.A1(_02530_),
    .A2(_02533_),
    .B1(_01591_),
    .Y(_02534_));
 sky130_fd_sc_hd__mux4_2 _07614_ (.A0(\rvsingle.dp.rf.rf[8][4] ),
    .A1(\rvsingle.dp.rf.rf[9][4] ),
    .A2(\rvsingle.dp.rf.rf[10][4] ),
    .A3(\rvsingle.dp.rf.rf[11][4] ),
    .S0(_01416_),
    .S1(_01708_),
    .X(_02535_));
 sky130_fd_sc_hd__or2_2 _07615_ (.A(_01419_),
    .B(\rvsingle.dp.rf.rf[12][4] ),
    .X(_02536_));
 sky130_fd_sc_hd__o211ai_2 _07616_ (.A1(\rvsingle.dp.rf.rf[13][4] ),
    .A2(_01440_),
    .B1(_01436_),
    .C1(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__or2_2 _07617_ (.A(_01690_),
    .B(\rvsingle.dp.rf.rf[14][4] ),
    .X(_02538_));
 sky130_fd_sc_hd__o211ai_2 _07618_ (.A1(_01687_),
    .A2(\rvsingle.dp.rf.rf[15][4] ),
    .B1(_01708_),
    .C1(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__a31oi_2 _07619_ (.A1(_02537_),
    .A2(_02539_),
    .A3(_02273_),
    .B1(_01217_),
    .Y(_02540_));
 sky130_fd_sc_hd__o21ai_2 _07620_ (.A1(_01711_),
    .A2(_02535_),
    .B1(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__mux4_2 _07621_ (.A0(\rvsingle.dp.rf.rf[4][4] ),
    .A1(\rvsingle.dp.rf.rf[5][4] ),
    .A2(\rvsingle.dp.rf.rf[6][4] ),
    .A3(\rvsingle.dp.rf.rf[7][4] ),
    .S0(_01416_),
    .S1(_01300_),
    .X(_02542_));
 sky130_fd_sc_hd__buf_1 _07622_ (.A(_01206_),
    .X(_02543_));
 sky130_fd_sc_hd__o21a_2 _07623_ (.A1(_01828_),
    .A2(\rvsingle.dp.rf.rf[2][4] ),
    .B1(_01299_),
    .X(_02544_));
 sky130_fd_sc_hd__o21ai_2 _07624_ (.A1(\rvsingle.dp.rf.rf[3][4] ),
    .A2(_02288_),
    .B1(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__or2_2 _07625_ (.A(_01690_),
    .B(\rvsingle.dp.rf.rf[0][4] ),
    .X(_02546_));
 sky130_fd_sc_hd__o211ai_2 _07626_ (.A1(\rvsingle.dp.rf.rf[1][4] ),
    .A2(_02271_),
    .B1(_02268_),
    .C1(_02546_),
    .Y(_02547_));
 sky130_fd_sc_hd__a31oi_2 _07627_ (.A1(_02543_),
    .A2(_02545_),
    .A3(_02547_),
    .B1(_01446_),
    .Y(_02548_));
 sky130_fd_sc_hd__o21ai_2 _07628_ (.A1(_01422_),
    .A2(_02542_),
    .B1(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__nand3_2 _07629_ (.A(_01315_),
    .B(_02541_),
    .C(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__or2_2 _07630_ (.A(_01419_),
    .B(\rvsingle.dp.rf.rf[28][4] ),
    .X(_02551_));
 sky130_fd_sc_hd__o211ai_2 _07631_ (.A1(\rvsingle.dp.rf.rf[29][4] ),
    .A2(_02275_),
    .B1(_01436_),
    .C1(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__o21a_2 _07632_ (.A1(_01725_),
    .A2(\rvsingle.dp.rf.rf[30][4] ),
    .B1(_01198_),
    .X(_02553_));
 sky130_fd_sc_hd__o21ai_2 _07633_ (.A1(\rvsingle.dp.rf.rf[31][4] ),
    .A2(_02288_),
    .B1(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__a31oi_2 _07634_ (.A1(_02552_),
    .A2(_02554_),
    .A3(_02273_),
    .B1(_01217_),
    .Y(_02555_));
 sky130_fd_sc_hd__or2_2 _07635_ (.A(_01191_),
    .B(\rvsingle.dp.rf.rf[24][4] ),
    .X(_02556_));
 sky130_fd_sc_hd__o211ai_2 _07636_ (.A1(\rvsingle.dp.rf.rf[25][4] ),
    .A2(_01295_),
    .B1(_01308_),
    .C1(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__o21a_2 _07637_ (.A1(_01903_),
    .A2(\rvsingle.dp.rf.rf[26][4] ),
    .B1(_01243_),
    .X(_02558_));
 sky130_fd_sc_hd__o21ai_2 _07638_ (.A1(\rvsingle.dp.rf.rf[27][4] ),
    .A2(_01901_),
    .B1(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand3_2 _07639_ (.A(_01721_),
    .B(_02557_),
    .C(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__a21oi_2 _07640_ (.A1(_02555_),
    .A2(_02560_),
    .B1(_01315_),
    .Y(_02561_));
 sky130_fd_sc_hd__mux4_2 _07641_ (.A0(\rvsingle.dp.rf.rf[16][4] ),
    .A1(\rvsingle.dp.rf.rf[17][4] ),
    .A2(\rvsingle.dp.rf.rf[18][4] ),
    .A3(\rvsingle.dp.rf.rf[19][4] ),
    .S0(_02176_),
    .S1(_02162_),
    .X(_02562_));
 sky130_fd_sc_hd__or2_2 _07642_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[20][4] ),
    .X(_02563_));
 sky130_fd_sc_hd__o211ai_2 _07643_ (.A1(\rvsingle.dp.rf.rf[21][4] ),
    .A2(_01827_),
    .B1(_01308_),
    .C1(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__or2_2 _07644_ (.A(_01419_),
    .B(\rvsingle.dp.rf.rf[22][4] ),
    .X(_02565_));
 sky130_fd_sc_hd__o211ai_2 _07645_ (.A1(_01440_),
    .A2(\rvsingle.dp.rf.rf[23][4] ),
    .B1(_01696_),
    .C1(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__a31oi_2 _07646_ (.A1(_02564_),
    .A2(_02566_),
    .A3(_02291_),
    .B1(_01446_),
    .Y(_02567_));
 sky130_fd_sc_hd__o21ai_2 _07647_ (.A1(_01711_),
    .A2(_02562_),
    .B1(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__nand2_2 _07648_ (.A(_02561_),
    .B(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hd__and3_2 _07649_ (.A(_01246_),
    .B(_02550_),
    .C(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__o21ai_2 _07650_ (.A1(Instr[11]),
    .A2(_01078_),
    .B1(_02531_),
    .Y(_02571_));
 sky130_fd_sc_hd__o221ai_2 _07651_ (.A1(_02473_),
    .A2(_02318_),
    .B1(_01537_),
    .B2(_02571_),
    .C1(_02530_),
    .Y(_02572_));
 sky130_fd_sc_hd__nand2_2 _07652_ (.A(_02570_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__nand2_2 _07653_ (.A(_02550_),
    .B(_02569_),
    .Y(_02574_));
 sky130_fd_sc_hd__o221a_2 _07654_ (.A1(_02473_),
    .A2(_02318_),
    .B1(_01537_),
    .B2(_02571_),
    .C1(_02530_),
    .X(_02575_));
 sky130_fd_sc_hd__o22ai_2 _07655_ (.A1(_02469_),
    .A2(_02574_),
    .B1(_02534_),
    .B2(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__o21a_2 _07656_ (.A1(_02534_),
    .A2(_02573_),
    .B1(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__or2_2 _07657_ (.A(_01690_),
    .B(\rvsingle.dp.rf.rf[4][5] ),
    .X(_02578_));
 sky130_fd_sc_hd__o211ai_2 _07658_ (.A1(\rvsingle.dp.rf.rf[5][5] ),
    .A2(_02271_),
    .B1(_02268_),
    .C1(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__o21a_2 _07659_ (.A1(_01191_),
    .A2(\rvsingle.dp.rf.rf[6][5] ),
    .B1(_01299_),
    .X(_02580_));
 sky130_fd_sc_hd__o21ai_2 _07660_ (.A1(\rvsingle.dp.rf.rf[7][5] ),
    .A2(_01440_),
    .B1(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__a31o_2 _07661_ (.A1(_02579_),
    .A2(_01444_),
    .A3(_02581_),
    .B1(_01215_),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_2 _07662_ (.A0(\rvsingle.dp.rf.rf[0][5] ),
    .A1(\rvsingle.dp.rf.rf[1][5] ),
    .S(_02176_),
    .X(_02583_));
 sky130_fd_sc_hd__or2_2 _07663_ (.A(_01419_),
    .B(\rvsingle.dp.rf.rf[2][5] ),
    .X(_02584_));
 sky130_fd_sc_hd__o211a_2 _07664_ (.A1(_01687_),
    .A2(\rvsingle.dp.rf.rf[3][5] ),
    .B1(_01455_),
    .C1(_02584_),
    .X(_02585_));
 sky130_fd_sc_hd__a211oi_2 _07665_ (.A1(_02583_),
    .A2(_01689_),
    .B1(_01702_),
    .C1(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__mux2_2 _07666_ (.A0(\rvsingle.dp.rf.rf[8][5] ),
    .A1(\rvsingle.dp.rf.rf[9][5] ),
    .S(_01426_),
    .X(_02587_));
 sky130_fd_sc_hd__or2_2 _07667_ (.A(_01349_),
    .B(\rvsingle.dp.rf.rf[10][5] ),
    .X(_02588_));
 sky130_fd_sc_hd__o211a_2 _07668_ (.A1(_02271_),
    .A2(\rvsingle.dp.rf.rf[11][5] ),
    .B1(_01300_),
    .C1(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__a211oi_2 _07669_ (.A1(_02587_),
    .A2(_01689_),
    .B1(_01702_),
    .C1(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__mux4_2 _07670_ (.A0(\rvsingle.dp.rf.rf[12][5] ),
    .A1(\rvsingle.dp.rf.rf[13][5] ),
    .A2(\rvsingle.dp.rf.rf[14][5] ),
    .A3(\rvsingle.dp.rf.rf[15][5] ),
    .S0(_01462_),
    .S1(_01727_),
    .X(_02591_));
 sky130_fd_sc_hd__o21ai_2 _07671_ (.A1(_01721_),
    .A2(_02591_),
    .B1(_02438_),
    .Y(_02592_));
 sky130_fd_sc_hd__o22ai_2 _07672_ (.A1(_02582_),
    .A2(_02586_),
    .B1(_02590_),
    .B2(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__mux4_2 _07673_ (.A0(\rvsingle.dp.rf.rf[24][5] ),
    .A1(\rvsingle.dp.rf.rf[25][5] ),
    .A2(\rvsingle.dp.rf.rf[26][5] ),
    .A3(\rvsingle.dp.rf.rf[27][5] ),
    .S0(_01328_),
    .S1(_01455_),
    .X(_02594_));
 sky130_fd_sc_hd__mux2_2 _07674_ (.A0(\rvsingle.dp.rf.rf[28][5] ),
    .A1(\rvsingle.dp.rf.rf[29][5] ),
    .S(_01419_),
    .X(_02595_));
 sky130_fd_sc_hd__or2_2 _07675_ (.A(_01327_),
    .B(\rvsingle.dp.rf.rf[30][5] ),
    .X(_02596_));
 sky130_fd_sc_hd__o211a_2 _07676_ (.A1(_01294_),
    .A2(\rvsingle.dp.rf.rf[31][5] ),
    .B1(_01243_),
    .C1(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__a211o_2 _07677_ (.A1(_02595_),
    .A2(_02285_),
    .B1(_01206_),
    .C1(_02597_),
    .X(_02598_));
 sky130_fd_sc_hd__o211ai_2 _07678_ (.A1(_02302_),
    .A2(_02594_),
    .B1(_02438_),
    .C1(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__mux4_2 _07679_ (.A0(\rvsingle.dp.rf.rf[20][5] ),
    .A1(\rvsingle.dp.rf.rf[21][5] ),
    .A2(\rvsingle.dp.rf.rf[22][5] ),
    .A3(\rvsingle.dp.rf.rf[23][5] ),
    .S0(_02450_),
    .S1(_01455_),
    .X(_02600_));
 sky130_fd_sc_hd__or2_2 _07680_ (.A(_01690_),
    .B(\rvsingle.dp.rf.rf[16][5] ),
    .X(_02601_));
 sky130_fd_sc_hd__o211ai_2 _07681_ (.A1(\rvsingle.dp.rf.rf[17][5] ),
    .A2(_02271_),
    .B1(_02268_),
    .C1(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__or2_2 _07682_ (.A(_01690_),
    .B(\rvsingle.dp.rf.rf[18][5] ),
    .X(_02603_));
 sky130_fd_sc_hd__o211ai_2 _07683_ (.A1(_01687_),
    .A2(\rvsingle.dp.rf.rf[19][5] ),
    .B1(_01455_),
    .C1(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__a31oi_2 _07684_ (.A1(_01460_),
    .A2(_02602_),
    .A3(_02604_),
    .B1(_01215_),
    .Y(_02605_));
 sky130_fd_sc_hd__o21ai_2 _07685_ (.A1(_01422_),
    .A2(_02600_),
    .B1(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__nand3_2 _07686_ (.A(_02599_),
    .B(_02606_),
    .C(_01187_),
    .Y(_02607_));
 sky130_fd_sc_hd__o21ai_2 _07687_ (.A1(_01450_),
    .A2(_02593_),
    .B1(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_2 _07688_ (.A(_02375_),
    .B(Instr[25]),
    .Y(_02609_));
 sky130_fd_sc_hd__nor2_2 _07689_ (.A(_01862_),
    .B(\rvsingle.dp.rf.rf[10][5] ),
    .Y(_02610_));
 sky130_fd_sc_hd__o21ai_2 _07690_ (.A1(\rvsingle.dp.rf.rf[11][5] ),
    .A2(_01087_),
    .B1(_01654_),
    .Y(_02611_));
 sky130_fd_sc_hd__or2b_2 _07691_ (.A(\rvsingle.dp.rf.rf[9][5] ),
    .B_N(_01752_),
    .X(_02612_));
 sky130_fd_sc_hd__o211ai_2 _07692_ (.A1(_01847_),
    .A2(\rvsingle.dp.rf.rf[8][5] ),
    .B1(_02612_),
    .C1(_01667_),
    .Y(_02613_));
 sky130_fd_sc_hd__o211ai_2 _07693_ (.A1(_02610_),
    .A2(_02611_),
    .B1(_02613_),
    .C1(_02329_),
    .Y(_02614_));
 sky130_fd_sc_hd__nor2_2 _07694_ (.A(_01125_),
    .B(\rvsingle.dp.rf.rf[14][5] ),
    .Y(_02615_));
 sky130_fd_sc_hd__and2b_2 _07695_ (.A_N(\rvsingle.dp.rf.rf[15][5] ),
    .B(_01779_),
    .X(_02616_));
 sky130_fd_sc_hd__o21ba_2 _07696_ (.A1(_01096_),
    .A2(\rvsingle.dp.rf.rf[12][5] ),
    .B1_N(_01103_),
    .X(_02617_));
 sky130_fd_sc_hd__o21ai_2 _07697_ (.A1(_01645_),
    .A2(\rvsingle.dp.rf.rf[13][5] ),
    .B1(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__o311ai_2 _07698_ (.A1(_01542_),
    .A2(_02615_),
    .A3(_02616_),
    .B1(_01502_),
    .C1(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__nand3_2 _07699_ (.A(_02614_),
    .B(_02491_),
    .C(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__o21a_2 _07700_ (.A1(_01566_),
    .A2(\rvsingle.dp.rf.rf[6][5] ),
    .B1(_01258_),
    .X(_02621_));
 sky130_fd_sc_hd__o21a_2 _07701_ (.A1(_02379_),
    .A2(\rvsingle.dp.rf.rf[7][5] ),
    .B1(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__o21bai_2 _07702_ (.A1(_01125_),
    .A2(\rvsingle.dp.rf.rf[4][5] ),
    .B1_N(_01519_),
    .Y(_02623_));
 sky130_fd_sc_hd__and2b_2 _07703_ (.A_N(\rvsingle.dp.rf.rf[5][5] ),
    .B(_01594_),
    .X(_02624_));
 sky130_fd_sc_hd__o21ai_2 _07704_ (.A1(_02623_),
    .A2(_02624_),
    .B1(_01111_),
    .Y(_02625_));
 sky130_fd_sc_hd__nor2_2 _07705_ (.A(_01797_),
    .B(\rvsingle.dp.rf.rf[0][5] ),
    .Y(_02626_));
 sky130_fd_sc_hd__buf_1 _07706_ (.A(_01135_),
    .X(_02627_));
 sky130_fd_sc_hd__and2b_2 _07707_ (.A_N(\rvsingle.dp.rf.rf[1][5] ),
    .B(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__or2b_2 _07708_ (.A(\rvsingle.dp.rf.rf[3][5] ),
    .B_N(_01606_),
    .X(_02629_));
 sky130_fd_sc_hd__o211ai_2 _07709_ (.A1(_01607_),
    .A2(\rvsingle.dp.rf.rf[2][5] ),
    .B1(_01596_),
    .C1(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__o311ai_2 _07710_ (.A1(_01520_),
    .A2(_02626_),
    .A3(_02628_),
    .B1(_01564_),
    .C1(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__o211ai_2 _07711_ (.A1(_02622_),
    .A2(_02625_),
    .B1(_02364_),
    .C1(_02631_),
    .Y(_02632_));
 sky130_fd_sc_hd__nand3_2 _07712_ (.A(_01377_),
    .B(_02620_),
    .C(_02632_),
    .Y(_02633_));
 sky130_fd_sc_hd__nor2_2 _07713_ (.A(_01862_),
    .B(\rvsingle.dp.rf.rf[30][5] ),
    .Y(_02634_));
 sky130_fd_sc_hd__o21ai_2 _07714_ (.A1(\rvsingle.dp.rf.rf[31][5] ),
    .A2(_01860_),
    .B1(_01880_),
    .Y(_02635_));
 sky130_fd_sc_hd__or2b_2 _07715_ (.A(\rvsingle.dp.rf.rf[29][5] ),
    .B_N(_01752_),
    .X(_02636_));
 sky130_fd_sc_hd__o211ai_2 _07716_ (.A1(_01675_),
    .A2(\rvsingle.dp.rf.rf[28][5] ),
    .B1(_02636_),
    .C1(_01667_),
    .Y(_02637_));
 sky130_fd_sc_hd__o211ai_2 _07717_ (.A1(_02634_),
    .A2(_02635_),
    .B1(_02637_),
    .C1(_02323_),
    .Y(_02638_));
 sky130_fd_sc_hd__nor2_2 _07718_ (.A(_01743_),
    .B(\rvsingle.dp.rf.rf[24][5] ),
    .Y(_02639_));
 sky130_fd_sc_hd__and2b_2 _07719_ (.A_N(\rvsingle.dp.rf.rf[25][5] ),
    .B(_01877_),
    .X(_02640_));
 sky130_fd_sc_hd__or2b_2 _07720_ (.A(\rvsingle.dp.rf.rf[27][5] ),
    .B_N(_01606_),
    .X(_02641_));
 sky130_fd_sc_hd__o211ai_2 _07721_ (.A1(_01797_),
    .A2(\rvsingle.dp.rf.rf[26][5] ),
    .B1(_01647_),
    .C1(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__o311ai_2 _07722_ (.A1(_02337_),
    .A2(_02639_),
    .A3(_02640_),
    .B1(_01564_),
    .C1(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand3_2 _07723_ (.A(_02638_),
    .B(_02643_),
    .C(_02491_),
    .Y(_02644_));
 sky130_fd_sc_hd__inv_2 _07724_ (.A(\rvsingle.dp.rf.rf[21][5] ),
    .Y(_02645_));
 sky130_fd_sc_hd__nor2_2 _07725_ (.A(_01607_),
    .B(\rvsingle.dp.rf.rf[20][5] ),
    .Y(_02646_));
 sky130_fd_sc_hd__a211oi_2 _07726_ (.A1(_02645_),
    .A2(_01780_),
    .B1(_02337_),
    .C1(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__o21ai_2 _07727_ (.A1(_01769_),
    .A2(\rvsingle.dp.rf.rf[22][5] ),
    .B1(_01104_),
    .Y(_02648_));
 sky130_fd_sc_hd__and2b_2 _07728_ (.A_N(\rvsingle.dp.rf.rf[23][5] ),
    .B(_02627_),
    .X(_02649_));
 sky130_fd_sc_hd__o21ai_2 _07729_ (.A1(_02648_),
    .A2(_02649_),
    .B1(_01502_),
    .Y(_02650_));
 sky130_fd_sc_hd__nor2_2 _07730_ (.A(_01650_),
    .B(\rvsingle.dp.rf.rf[16][5] ),
    .Y(_02651_));
 sky130_fd_sc_hd__and2b_2 _07731_ (.A_N(\rvsingle.dp.rf.rf[17][5] ),
    .B(_01566_),
    .X(_02652_));
 sky130_fd_sc_hd__o21a_2 _07732_ (.A1(_01752_),
    .A2(\rvsingle.dp.rf.rf[18][5] ),
    .B1(_01610_),
    .X(_02653_));
 sky130_fd_sc_hd__o21ai_2 _07733_ (.A1(\rvsingle.dp.rf.rf[19][5] ),
    .A2(_01087_),
    .B1(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__o311ai_2 _07734_ (.A1(_01777_),
    .A2(_02651_),
    .A3(_02652_),
    .B1(_01599_),
    .C1(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__o211ai_2 _07735_ (.A1(_02647_),
    .A2(_02650_),
    .B1(_02364_),
    .C1(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand3_2 _07736_ (.A(_02644_),
    .B(_02656_),
    .C(_01145_),
    .Y(_02657_));
 sky130_fd_sc_hd__nand4_2 _07737_ (.A(_02633_),
    .B(_01083_),
    .C(_02505_),
    .D(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__o211a_2 _07738_ (.A1(_01065_),
    .A2(_01074_),
    .B1(_02609_),
    .C1(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__a21oi_2 _07739_ (.A1(_02609_),
    .A2(_02658_),
    .B1(_01591_),
    .Y(_02660_));
 sky130_fd_sc_hd__o22ai_2 _07740_ (.A1(_02469_),
    .A2(_02608_),
    .B1(_02659_),
    .B2(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__o211ai_2 _07741_ (.A1(_01150_),
    .A2(_01139_),
    .B1(_02657_),
    .C1(_02633_),
    .Y(_02662_));
 sky130_fd_sc_hd__nand2_2 _07742_ (.A(_02662_),
    .B(_01481_),
    .Y(_02663_));
 sky130_fd_sc_hd__o211ai_2 _07743_ (.A1(Instr[25]),
    .A2(_01537_),
    .B1(_01183_),
    .C1(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hd__o211a_2 _07744_ (.A1(_02315_),
    .A2(_02593_),
    .B1(_02607_),
    .C1(_01246_),
    .X(_02665_));
 sky130_fd_sc_hd__o221ai_2 _07745_ (.A1(_01065_),
    .A2(_01074_),
    .B1(_01178_),
    .B2(_02662_),
    .C1(_02609_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand3_2 _07746_ (.A(_02664_),
    .B(_02665_),
    .C(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand4_2 _07747_ (.A(_02476_),
    .B(_02577_),
    .C(_02661_),
    .D(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__mux2_2 _07748_ (.A0(\rvsingle.dp.rf.rf[0][3] ),
    .A1(\rvsingle.dp.rf.rf[1][3] ),
    .S(_01241_),
    .X(_02669_));
 sky130_fd_sc_hd__or2_2 _07749_ (.A(_01828_),
    .B(\rvsingle.dp.rf.rf[2][3] ),
    .X(_02670_));
 sky130_fd_sc_hd__o211a_2 _07750_ (.A1(_02288_),
    .A2(\rvsingle.dp.rf.rf[3][3] ),
    .B1(_01433_),
    .C1(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__a211oi_2 _07751_ (.A1(_02669_),
    .A2(_01437_),
    .B1(_01229_),
    .C1(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__mux4_2 _07752_ (.A0(\rvsingle.dp.rf.rf[4][3] ),
    .A1(\rvsingle.dp.rf.rf[5][3] ),
    .A2(\rvsingle.dp.rf.rf[6][3] ),
    .A3(\rvsingle.dp.rf.rf[7][3] ),
    .S0(_01903_),
    .S1(_01470_),
    .X(_02673_));
 sky130_fd_sc_hd__o21ai_2 _07753_ (.A1(_01207_),
    .A2(_02673_),
    .B1(_02447_),
    .Y(_02674_));
 sky130_fd_sc_hd__mux4_2 _07754_ (.A0(\rvsingle.dp.rf.rf[8][3] ),
    .A1(\rvsingle.dp.rf.rf[9][3] ),
    .A2(\rvsingle.dp.rf.rf[10][3] ),
    .A3(\rvsingle.dp.rf.rf[11][3] ),
    .S0(_02176_),
    .S1(_01696_),
    .X(_02675_));
 sky130_fd_sc_hd__or2_2 _07755_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[12][3] ),
    .X(_02676_));
 sky130_fd_sc_hd__o211ai_2 _07756_ (.A1(\rvsingle.dp.rf.rf[13][3] ),
    .A2(_02288_),
    .B1(_01436_),
    .C1(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__or2_2 _07757_ (.A(_01419_),
    .B(\rvsingle.dp.rf.rf[14][3] ),
    .X(_02678_));
 sky130_fd_sc_hd__o211ai_2 _07758_ (.A1(_02271_),
    .A2(\rvsingle.dp.rf.rf[15][3] ),
    .B1(_01300_),
    .C1(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__a31oi_2 _07759_ (.A1(_02677_),
    .A2(_02679_),
    .A3(_02291_),
    .B1(_01217_),
    .Y(_02680_));
 sky130_fd_sc_hd__o21ai_2 _07760_ (.A1(_01711_),
    .A2(_02675_),
    .B1(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__o21ai_2 _07761_ (.A1(_02672_),
    .A2(_02674_),
    .B1(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__mux2_2 _07762_ (.A0(\rvsingle.dp.rf.rf[20][3] ),
    .A1(\rvsingle.dp.rf.rf[21][3] ),
    .S(_01335_),
    .X(_02683_));
 sky130_fd_sc_hd__or2_2 _07763_ (.A(_01828_),
    .B(\rvsingle.dp.rf.rf[22][3] ),
    .X(_02684_));
 sky130_fd_sc_hd__o211a_2 _07764_ (.A1(_01827_),
    .A2(\rvsingle.dp.rf.rf[23][3] ),
    .B1(_01808_),
    .C1(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__a211oi_2 _07765_ (.A1(_02683_),
    .A2(_01437_),
    .B1(_01721_),
    .C1(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__mux4_2 _07766_ (.A0(\rvsingle.dp.rf.rf[16][3] ),
    .A1(\rvsingle.dp.rf.rf[17][3] ),
    .A2(\rvsingle.dp.rf.rf[18][3] ),
    .A3(\rvsingle.dp.rf.rf[19][3] ),
    .S0(_01328_),
    .S1(_01455_),
    .X(_02687_));
 sky130_fd_sc_hd__o21ai_2 _07767_ (.A1(_02302_),
    .A2(_02687_),
    .B1(_02447_),
    .Y(_02688_));
 sky130_fd_sc_hd__mux4_2 _07768_ (.A0(\rvsingle.dp.rf.rf[24][3] ),
    .A1(\rvsingle.dp.rf.rf[25][3] ),
    .A2(\rvsingle.dp.rf.rf[26][3] ),
    .A3(\rvsingle.dp.rf.rf[27][3] ),
    .S0(_02450_),
    .S1(_01708_),
    .X(_02689_));
 sky130_fd_sc_hd__mux2_2 _07769_ (.A0(\rvsingle.dp.rf.rf[28][3] ),
    .A1(\rvsingle.dp.rf.rf[29][3] ),
    .S(_01419_),
    .X(_02690_));
 sky130_fd_sc_hd__o21a_2 _07770_ (.A1(_01425_),
    .A2(\rvsingle.dp.rf.rf[30][3] ),
    .B1(_01197_),
    .X(_02691_));
 sky130_fd_sc_hd__o21a_2 _07771_ (.A1(_01423_),
    .A2(\rvsingle.dp.rf.rf[31][3] ),
    .B1(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__a211o_2 _07772_ (.A1(_02690_),
    .A2(_02285_),
    .B1(_01206_),
    .C1(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__o211ai_2 _07773_ (.A1(_02302_),
    .A2(_02689_),
    .B1(_02693_),
    .C1(_02438_),
    .Y(_02694_));
 sky130_fd_sc_hd__o211ai_2 _07774_ (.A1(_02686_),
    .A2(_02688_),
    .B1(_01187_),
    .C1(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__o21ai_2 _07775_ (.A1(_01188_),
    .A2(_02682_),
    .B1(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hd__a31o_2 _07776_ (.A1(_01076_),
    .A2(_01071_),
    .A3(_01062_),
    .B1(_01115_),
    .X(_02697_));
 sky130_fd_sc_hd__o21ai_2 _07777_ (.A1(Instr[10]),
    .A2(_01078_),
    .B1(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__nor2_2 _07778_ (.A(_01097_),
    .B(\rvsingle.dp.rf.rf[8][3] ),
    .Y(_02699_));
 sky130_fd_sc_hd__o21ai_2 _07779_ (.A1(\rvsingle.dp.rf.rf[9][3] ),
    .A2(_01087_),
    .B1(_01667_),
    .Y(_02700_));
 sky130_fd_sc_hd__or2_2 _07780_ (.A(_01752_),
    .B(\rvsingle.dp.rf.rf[10][3] ),
    .X(_02701_));
 sky130_fd_sc_hd__o211ai_2 _07781_ (.A1(_01087_),
    .A2(\rvsingle.dp.rf.rf[11][3] ),
    .B1(_01611_),
    .C1(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__o211ai_2 _07782_ (.A1(_02699_),
    .A2(_02700_),
    .B1(_01564_),
    .C1(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__and2b_2 _07783_ (.A_N(\rvsingle.dp.rf.rf[15][3] ),
    .B(_01566_),
    .X(_02704_));
 sky130_fd_sc_hd__o21ai_2 _07784_ (.A1(_01650_),
    .A2(\rvsingle.dp.rf.rf[14][3] ),
    .B1(_01647_),
    .Y(_02705_));
 sky130_fd_sc_hd__nor2_2 _07785_ (.A(_01607_),
    .B(\rvsingle.dp.rf.rf[12][3] ),
    .Y(_02706_));
 sky130_fd_sc_hd__o21ai_2 _07786_ (.A1(\rvsingle.dp.rf.rf[13][3] ),
    .A2(_01645_),
    .B1(_01667_),
    .Y(_02707_));
 sky130_fd_sc_hd__o221ai_2 _07787_ (.A1(_02704_),
    .A2(_02705_),
    .B1(_02706_),
    .B2(_02707_),
    .C1(_01111_),
    .Y(_02708_));
 sky130_fd_sc_hd__nand3_2 _07788_ (.A(_02703_),
    .B(_02491_),
    .C(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__nor2_2 _07789_ (.A(_02005_),
    .B(\rvsingle.dp.rf.rf[0][3] ),
    .Y(_02710_));
 sky130_fd_sc_hd__and2b_2 _07790_ (.A_N(\rvsingle.dp.rf.rf[1][3] ),
    .B(_01566_),
    .X(_02711_));
 sky130_fd_sc_hd__or2b_2 _07791_ (.A(\rvsingle.dp.rf.rf[3][3] ),
    .B_N(_01606_),
    .X(_02712_));
 sky130_fd_sc_hd__o211ai_2 _07792_ (.A1(_01125_),
    .A2(\rvsingle.dp.rf.rf[2][3] ),
    .B1(_01647_),
    .C1(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__o311ai_2 _07793_ (.A1(_02031_),
    .A2(_02710_),
    .A3(_02711_),
    .B1(_01599_),
    .C1(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__nor2_2 _07794_ (.A(_01125_),
    .B(\rvsingle.dp.rf.rf[4][3] ),
    .Y(_02715_));
 sky130_fd_sc_hd__and2b_2 _07795_ (.A_N(\rvsingle.dp.rf.rf[5][3] ),
    .B(_01779_),
    .X(_02716_));
 sky130_fd_sc_hd__or2b_2 _07796_ (.A(\rvsingle.dp.rf.rf[7][3] ),
    .B_N(_01606_),
    .X(_02717_));
 sky130_fd_sc_hd__o211ai_2 _07797_ (.A1(_01743_),
    .A2(\rvsingle.dp.rf.rf[6][3] ),
    .B1(_01647_),
    .C1(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__o311ai_2 _07798_ (.A1(_02031_),
    .A2(_02715_),
    .A3(_02716_),
    .B1(_01502_),
    .C1(_02718_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand3_2 _07799_ (.A(_02364_),
    .B(_02714_),
    .C(_02719_),
    .Y(_02720_));
 sky130_fd_sc_hd__nand3_2 _07800_ (.A(_01376_),
    .B(_02709_),
    .C(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__nor2_2 _07801_ (.A(_01642_),
    .B(\rvsingle.dp.rf.rf[28][3] ),
    .Y(_02722_));
 sky130_fd_sc_hd__and2b_2 _07802_ (.A_N(\rvsingle.dp.rf.rf[29][3] ),
    .B(_01498_),
    .X(_02723_));
 sky130_fd_sc_hd__or2b_2 _07803_ (.A(\rvsingle.dp.rf.rf[31][3] ),
    .B_N(_01752_),
    .X(_02724_));
 sky130_fd_sc_hd__o211ai_2 _07804_ (.A1(_01753_),
    .A2(\rvsingle.dp.rf.rf[30][3] ),
    .B1(_01596_),
    .C1(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__o311ai_2 _07805_ (.A1(_01520_),
    .A2(_02722_),
    .A3(_02723_),
    .B1(_01111_),
    .C1(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__nor2_2 _07806_ (.A(_01125_),
    .B(\rvsingle.dp.rf.rf[24][3] ),
    .Y(_02727_));
 sky130_fd_sc_hd__and2b_2 _07807_ (.A_N(\rvsingle.dp.rf.rf[25][3] ),
    .B(_01779_),
    .X(_02728_));
 sky130_fd_sc_hd__or2b_2 _07808_ (.A(\rvsingle.dp.rf.rf[27][3] ),
    .B_N(_01606_),
    .X(_02729_));
 sky130_fd_sc_hd__o211ai_2 _07809_ (.A1(_01797_),
    .A2(\rvsingle.dp.rf.rf[26][3] ),
    .B1(_01647_),
    .C1(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__o311ai_2 _07810_ (.A1(_02337_),
    .A2(_02727_),
    .A3(_02728_),
    .B1(_01599_),
    .C1(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__nand3_2 _07811_ (.A(_02726_),
    .B(_02731_),
    .C(_02491_),
    .Y(_02732_));
 sky130_fd_sc_hd__inv_2 _07812_ (.A(\rvsingle.dp.rf.rf[23][3] ),
    .Y(_02733_));
 sky130_fd_sc_hd__nor2_2 _07813_ (.A(_01797_),
    .B(\rvsingle.dp.rf.rf[22][3] ),
    .Y(_02734_));
 sky130_fd_sc_hd__a211oi_2 _07814_ (.A1(_02733_),
    .A2(_02030_),
    .B1(_01542_),
    .C1(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__o21bai_2 _07815_ (.A1(_01602_),
    .A2(\rvsingle.dp.rf.rf[20][3] ),
    .B1_N(_01258_),
    .Y(_02736_));
 sky130_fd_sc_hd__and2b_2 _07816_ (.A_N(\rvsingle.dp.rf.rf[21][3] ),
    .B(_02627_),
    .X(_02737_));
 sky130_fd_sc_hd__o21ai_2 _07817_ (.A1(_02736_),
    .A2(_02737_),
    .B1(_01502_),
    .Y(_02738_));
 sky130_fd_sc_hd__nor2_2 _07818_ (.A(_01650_),
    .B(\rvsingle.dp.rf.rf[16][3] ),
    .Y(_02739_));
 sky130_fd_sc_hd__and2b_2 _07819_ (.A_N(\rvsingle.dp.rf.rf[17][3] ),
    .B(_01544_),
    .X(_02740_));
 sky130_fd_sc_hd__or2b_2 _07820_ (.A(\rvsingle.dp.rf.rf[19][3] ),
    .B_N(_01124_),
    .X(_02741_));
 sky130_fd_sc_hd__o211ai_2 _07821_ (.A1(_01650_),
    .A2(\rvsingle.dp.rf.rf[18][3] ),
    .B1(_01104_),
    .C1(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__o311ai_2 _07822_ (.A1(_01777_),
    .A2(_02739_),
    .A3(_02740_),
    .B1(_01599_),
    .C1(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__o211ai_2 _07823_ (.A1(_02735_),
    .A2(_02738_),
    .B1(_02364_),
    .C1(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__nand3_2 _07824_ (.A(_02732_),
    .B(_02744_),
    .C(_01145_),
    .Y(_02745_));
 sky130_fd_sc_hd__nand4_2 _07825_ (.A(_02721_),
    .B(_01082_),
    .C(_01152_),
    .D(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__o221a_2 _07826_ (.A1(_01065_),
    .A2(_01074_),
    .B1(_01481_),
    .B2(_02698_),
    .C1(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__o21a_2 _07827_ (.A1(Instr[10]),
    .A2(_01078_),
    .B1(_02697_),
    .X(_02748_));
 sky130_fd_sc_hd__nand2_2 _07828_ (.A(_02375_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__a21oi_2 _07829_ (.A1(_02749_),
    .A2(_02746_),
    .B1(_01485_),
    .Y(_02750_));
 sky130_fd_sc_hd__o22ai_2 _07830_ (.A1(_02469_),
    .A2(_02696_),
    .B1(_02747_),
    .B2(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__nor2_2 _07831_ (.A(_02030_),
    .B(\rvsingle.dp.rf.rf[10][2] ),
    .Y(_02752_));
 sky130_fd_sc_hd__o21ai_2 _07832_ (.A1(\rvsingle.dp.rf.rf[11][2] ),
    .A2(_01539_),
    .B1(_02337_),
    .Y(_02753_));
 sky130_fd_sc_hd__or2_2 _07833_ (.A(_01381_),
    .B(\rvsingle.dp.rf.rf[8][2] ),
    .X(_02754_));
 sky130_fd_sc_hd__o211ai_2 _07834_ (.A1(\rvsingle.dp.rf.rf[9][2] ),
    .A2(_01539_),
    .B1(_01542_),
    .C1(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__o211ai_2 _07835_ (.A1(_02752_),
    .A2(_02753_),
    .B1(_01131_),
    .C1(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__o21ba_2 _07836_ (.A1(_01594_),
    .A2(\rvsingle.dp.rf.rf[12][2] ),
    .B1_N(_01258_),
    .X(_02757_));
 sky130_fd_sc_hd__o21ai_2 _07837_ (.A1(_01508_),
    .A2(\rvsingle.dp.rf.rf[13][2] ),
    .B1(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__o21a_2 _07838_ (.A1(_02627_),
    .A2(\rvsingle.dp.rf.rf[14][2] ),
    .B1(_01519_),
    .X(_02759_));
 sky130_fd_sc_hd__o21ai_2 _07839_ (.A1(\rvsingle.dp.rf.rf[15][2] ),
    .A2(_01539_),
    .B1(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__nand3_2 _07840_ (.A(_02758_),
    .B(_02410_),
    .C(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__nand3_2 _07841_ (.A(_02756_),
    .B(_01505_),
    .C(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__o21bai_2 _07842_ (.A1(_01607_),
    .A2(\rvsingle.dp.rf.rf[0][2] ),
    .B1_N(_01489_),
    .Y(_02763_));
 sky130_fd_sc_hd__and2b_2 _07843_ (.A_N(\rvsingle.dp.rf.rf[1][2] ),
    .B(_01613_),
    .X(_02764_));
 sky130_fd_sc_hd__o21ai_2 _07844_ (.A1(_02763_),
    .A2(_02764_),
    .B1(_02329_),
    .Y(_02765_));
 sky130_fd_sc_hd__or2b_2 _07845_ (.A(\rvsingle.dp.rf.rf[3][2] ),
    .B_N(_02627_),
    .X(_02766_));
 sky130_fd_sc_hd__o211a_2 _07846_ (.A1(_01567_),
    .A2(\rvsingle.dp.rf.rf[2][2] ),
    .B1(_02031_),
    .C1(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_2 _07847_ (.A(_01675_),
    .B(\rvsingle.dp.rf.rf[4][2] ),
    .Y(_02768_));
 sky130_fd_sc_hd__and2b_2 _07848_ (.A_N(\rvsingle.dp.rf.rf[5][2] ),
    .B(_01492_),
    .X(_02769_));
 sky130_fd_sc_hd__or2b_2 _07849_ (.A(\rvsingle.dp.rf.rf[7][2] ),
    .B_N(_01096_),
    .X(_02770_));
 sky130_fd_sc_hd__o211ai_2 _07850_ (.A1(_01148_),
    .A2(\rvsingle.dp.rf.rf[6][2] ),
    .B1(_01611_),
    .C1(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__o311ai_2 _07851_ (.A1(_01490_),
    .A2(_02768_),
    .A3(_02769_),
    .B1(_01111_),
    .C1(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__o211ai_2 _07852_ (.A1(_02765_),
    .A2(_02767_),
    .B1(_02364_),
    .C1(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__nand3_2 _07853_ (.A(_01377_),
    .B(_02762_),
    .C(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__nor2_2 _07854_ (.A(_01499_),
    .B(\rvsingle.dp.rf.rf[30][2] ),
    .Y(_02775_));
 sky130_fd_sc_hd__o21ai_2 _07855_ (.A1(\rvsingle.dp.rf.rf[31][2] ),
    .A2(_01539_),
    .B1(_01520_),
    .Y(_02776_));
 sky130_fd_sc_hd__or2_2 _07856_ (.A(_01877_),
    .B(\rvsingle.dp.rf.rf[28][2] ),
    .X(_02777_));
 sky130_fd_sc_hd__o211ai_2 _07857_ (.A1(\rvsingle.dp.rf.rf[29][2] ),
    .A2(_01508_),
    .B1(_02395_),
    .C1(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__o211ai_2 _07858_ (.A1(_02775_),
    .A2(_02776_),
    .B1(_02410_),
    .C1(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__nor2_2 _07859_ (.A(_01097_),
    .B(\rvsingle.dp.rf.rf[24][2] ),
    .Y(_02780_));
 sky130_fd_sc_hd__and2b_2 _07860_ (.A_N(\rvsingle.dp.rf.rf[25][2] ),
    .B(_01613_),
    .X(_02781_));
 sky130_fd_sc_hd__or2b_2 _07861_ (.A(\rvsingle.dp.rf.rf[27][2] ),
    .B_N(_01381_),
    .X(_02782_));
 sky130_fd_sc_hd__o211ai_2 _07862_ (.A1(_01862_),
    .A2(\rvsingle.dp.rf.rf[26][2] ),
    .B1(_01880_),
    .C1(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__o311ai_2 _07863_ (.A1(_01552_),
    .A2(_02780_),
    .A3(_02781_),
    .B1(_02329_),
    .C1(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__nand3_2 _07864_ (.A(_02779_),
    .B(_02784_),
    .C(_01505_),
    .Y(_02785_));
 sky130_fd_sc_hd__nor2_2 _07865_ (.A(_01847_),
    .B(\rvsingle.dp.rf.rf[16][2] ),
    .Y(_02786_));
 sky130_fd_sc_hd__and2b_2 _07866_ (.A_N(\rvsingle.dp.rf.rf[17][2] ),
    .B(_01594_),
    .X(_02787_));
 sky130_fd_sc_hd__or2b_2 _07867_ (.A(\rvsingle.dp.rf.rf[19][2] ),
    .B_N(_01096_),
    .X(_02788_));
 sky130_fd_sc_hd__o211ai_2 _07868_ (.A1(_01148_),
    .A2(\rvsingle.dp.rf.rf[18][2] ),
    .B1(_01611_),
    .C1(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__o311ai_2 _07869_ (.A1(_01490_),
    .A2(_02786_),
    .A3(_02787_),
    .B1(_02329_),
    .C1(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__or2b_2 _07870_ (.A(\rvsingle.dp.rf.rf[21][2] ),
    .B_N(_01544_),
    .X(_02791_));
 sky130_fd_sc_hd__o211ai_2 _07871_ (.A1(_01567_),
    .A2(\rvsingle.dp.rf.rf[20][2] ),
    .B1(_02791_),
    .C1(_02395_),
    .Y(_02792_));
 sky130_fd_sc_hd__or2b_2 _07872_ (.A(\rvsingle.dp.rf.rf[23][2] ),
    .B_N(_01544_),
    .X(_02793_));
 sky130_fd_sc_hd__o211ai_2 _07873_ (.A1(_01558_),
    .A2(\rvsingle.dp.rf.rf[22][2] ),
    .B1(_01259_),
    .C1(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__nand3_2 _07874_ (.A(_02792_),
    .B(_02410_),
    .C(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__nand3_2 _07875_ (.A(_01156_),
    .B(_02790_),
    .C(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hd__nand3_2 _07876_ (.A(_02785_),
    .B(_02796_),
    .C(_01146_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand4_2 _07877_ (.A(_01152_),
    .B(_02774_),
    .C(_02797_),
    .D(_01082_),
    .Y(_02798_));
 sky130_fd_sc_hd__buf_1 _07878_ (.A(_01068_),
    .X(_02799_));
 sky130_fd_sc_hd__or4_2 _07879_ (.A(Instr[3]),
    .B(Instr[2]),
    .C(Instr[9]),
    .D(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__o21a_2 _07880_ (.A1(_01512_),
    .A2(_01069_),
    .B1(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__nand2_2 _07881_ (.A(_02801_),
    .B(_02375_),
    .Y(_02802_));
 sky130_fd_sc_hd__a21oi_2 _07882_ (.A1(_02798_),
    .A2(_02802_),
    .B1(_01485_),
    .Y(_02803_));
 sky130_fd_sc_hd__or2_2 _07883_ (.A(_01419_),
    .B(\rvsingle.dp.rf.rf[12][2] ),
    .X(_02804_));
 sky130_fd_sc_hd__o211ai_2 _07884_ (.A1(\rvsingle.dp.rf.rf[13][2] ),
    .A2(_01440_),
    .B1(_02268_),
    .C1(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__o21a_2 _07885_ (.A1(_01828_),
    .A2(\rvsingle.dp.rf.rf[14][2] ),
    .B1(_01299_),
    .X(_02806_));
 sky130_fd_sc_hd__o21ai_2 _07886_ (.A1(\rvsingle.dp.rf.rf[15][2] ),
    .A2(_02275_),
    .B1(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__a31oi_2 _07887_ (.A1(_02805_),
    .A2(_02273_),
    .A3(_02807_),
    .B1(_01217_),
    .Y(_02808_));
 sky130_fd_sc_hd__nor2_2 _07888_ (.A(_01726_),
    .B(\rvsingle.dp.rf.rf[8][2] ),
    .Y(_02809_));
 sky130_fd_sc_hd__o21ai_2 _07889_ (.A1(\rvsingle.dp.rf.rf[9][2] ),
    .A2(_02288_),
    .B1(_01308_),
    .Y(_02810_));
 sky130_fd_sc_hd__o21a_2 _07890_ (.A1(_01903_),
    .A2(\rvsingle.dp.rf.rf[10][2] ),
    .B1(_01243_),
    .X(_02811_));
 sky130_fd_sc_hd__o21ai_2 _07891_ (.A1(\rvsingle.dp.rf.rf[11][2] ),
    .A2(_01901_),
    .B1(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__o211ai_2 _07892_ (.A1(_02809_),
    .A2(_02810_),
    .B1(_02543_),
    .C1(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__nand2_2 _07893_ (.A(_02808_),
    .B(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__nor2_2 _07894_ (.A(_01420_),
    .B(\rvsingle.dp.rf.rf[2][2] ),
    .Y(_02815_));
 sky130_fd_sc_hd__o21ai_2 _07895_ (.A1(\rvsingle.dp.rf.rf[3][2] ),
    .A2(_02271_),
    .B1(_01300_),
    .Y(_02816_));
 sky130_fd_sc_hd__o21ba_2 _07896_ (.A1(_01725_),
    .A2(\rvsingle.dp.rf.rf[0][2] ),
    .B1_N(_01454_),
    .X(_02817_));
 sky130_fd_sc_hd__o21ai_2 _07897_ (.A1(_02275_),
    .A2(\rvsingle.dp.rf.rf[1][2] ),
    .B1(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__o21ai_2 _07898_ (.A1(_02815_),
    .A2(_02816_),
    .B1(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__nor2_2 _07899_ (.A(_01691_),
    .B(\rvsingle.dp.rf.rf[6][2] ),
    .Y(_02820_));
 sky130_fd_sc_hd__o21ai_2 _07900_ (.A1(\rvsingle.dp.rf.rf[7][2] ),
    .A2(_01687_),
    .B1(_01470_),
    .Y(_02821_));
 sky130_fd_sc_hd__nor2_2 _07901_ (.A(_01707_),
    .B(\rvsingle.dp.rf.rf[4][2] ),
    .Y(_02822_));
 sky130_fd_sc_hd__o21ai_2 _07902_ (.A1(\rvsingle.dp.rf.rf[5][2] ),
    .A2(_01687_),
    .B1(_02268_),
    .Y(_02823_));
 sky130_fd_sc_hd__o221ai_2 _07903_ (.A1(_02820_),
    .A2(_02821_),
    .B1(_02822_),
    .B2(_02823_),
    .C1(_01444_),
    .Y(_02824_));
 sky130_fd_sc_hd__o211ai_2 _07904_ (.A1(_01229_),
    .A2(_02819_),
    .B1(_02824_),
    .C1(_01217_),
    .Y(_02825_));
 sky130_fd_sc_hd__nand3_2 _07905_ (.A(_01315_),
    .B(_02814_),
    .C(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__nor2_2 _07906_ (.A(_01420_),
    .B(\rvsingle.dp.rf.rf[22][2] ),
    .Y(_02827_));
 sky130_fd_sc_hd__nor2_2 _07907_ (.A(\rvsingle.dp.rf.rf[23][2] ),
    .B(_01295_),
    .Y(_02828_));
 sky130_fd_sc_hd__or2_2 _07908_ (.A(_01349_),
    .B(\rvsingle.dp.rf.rf[20][2] ),
    .X(_02829_));
 sky130_fd_sc_hd__o211ai_2 _07909_ (.A1(\rvsingle.dp.rf.rf[21][2] ),
    .A2(_02275_),
    .B1(_01436_),
    .C1(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__o311a_2 _07910_ (.A1(_02827_),
    .A2(_01716_),
    .A3(_02828_),
    .B1(_02830_),
    .C1(_02291_),
    .X(_02831_));
 sky130_fd_sc_hd__or2b_2 _07911_ (.A(\rvsingle.dp.rf.rf[19][2] ),
    .B_N(_01191_),
    .X(_02832_));
 sky130_fd_sc_hd__o211ai_2 _07912_ (.A1(_01420_),
    .A2(\rvsingle.dp.rf.rf[18][2] ),
    .B1(_01696_),
    .C1(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__o21ba_2 _07913_ (.A1(_01462_),
    .A2(\rvsingle.dp.rf.rf[16][2] ),
    .B1_N(_01299_),
    .X(_02834_));
 sky130_fd_sc_hd__o21ai_2 _07914_ (.A1(_01827_),
    .A2(\rvsingle.dp.rf.rf[17][2] ),
    .B1(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__a31o_2 _07915_ (.A1(_02543_),
    .A2(_02833_),
    .A3(_02835_),
    .B1(_01215_),
    .X(_02836_));
 sky130_fd_sc_hd__o21ba_2 _07916_ (.A1(_01462_),
    .A2(\rvsingle.dp.rf.rf[24][2] ),
    .B1_N(_01299_),
    .X(_02837_));
 sky130_fd_sc_hd__o21a_2 _07917_ (.A1(_02303_),
    .A2(\rvsingle.dp.rf.rf[25][2] ),
    .B1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__or2_2 _07918_ (.A(_01191_),
    .B(\rvsingle.dp.rf.rf[26][2] ),
    .X(_02839_));
 sky130_fd_sc_hd__o211a_2 _07919_ (.A1(_02275_),
    .A2(\rvsingle.dp.rf.rf[27][2] ),
    .B1(_02162_),
    .C1(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__or2_2 _07920_ (.A(_01690_),
    .B(\rvsingle.dp.rf.rf[28][2] ),
    .X(_02841_));
 sky130_fd_sc_hd__o211ai_2 _07921_ (.A1(\rvsingle.dp.rf.rf[29][2] ),
    .A2(_01687_),
    .B1(_02268_),
    .C1(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__or2b_2 _07922_ (.A(\rvsingle.dp.rf.rf[31][2] ),
    .B_N(_01690_),
    .X(_02843_));
 sky130_fd_sc_hd__o211ai_2 _07923_ (.A1(_01335_),
    .A2(\rvsingle.dp.rf.rf[30][2] ),
    .B1(_01727_),
    .C1(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__a31oi_2 _07924_ (.A1(_02842_),
    .A2(_02844_),
    .A3(_01444_),
    .B1(_01216_),
    .Y(_02845_));
 sky130_fd_sc_hd__o31ai_2 _07925_ (.A1(_01702_),
    .A2(_02838_),
    .A3(_02840_),
    .B1(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__o211ai_2 _07926_ (.A1(_02831_),
    .A2(_02836_),
    .B1(_01187_),
    .C1(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__and3_2 _07927_ (.A(_01246_),
    .B(_02826_),
    .C(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__o21ai_2 _07928_ (.A1(_01113_),
    .A2(_01069_),
    .B1(_02800_),
    .Y(_02849_));
 sky130_fd_sc_hd__o211ai_2 _07929_ (.A1(_02849_),
    .A2(_01537_),
    .B1(_01591_),
    .C1(_02798_),
    .Y(_02850_));
 sky130_fd_sc_hd__nand2_2 _07930_ (.A(_02848_),
    .B(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__o21ai_2 _07931_ (.A1(_01870_),
    .A2(_02698_),
    .B1(_02746_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand2_2 _07932_ (.A(_02852_),
    .B(_01584_),
    .Y(_02853_));
 sky130_fd_sc_hd__o211a_2 _07933_ (.A1(_01188_),
    .A2(_02682_),
    .B1(_02695_),
    .C1(_01247_),
    .X(_02854_));
 sky130_fd_sc_hd__o221ai_2 _07934_ (.A1(_02473_),
    .A2(_02318_),
    .B1(_01537_),
    .B2(_02698_),
    .C1(_02746_),
    .Y(_02855_));
 sky130_fd_sc_hd__nand3_2 _07935_ (.A(_02853_),
    .B(_02854_),
    .C(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__o21ai_2 _07936_ (.A1(_02803_),
    .A2(_02851_),
    .B1(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__inv_2 _07937_ (.A(_02847_),
    .Y(_02858_));
 sky130_fd_sc_hd__a31o_2 _07938_ (.A1(_01316_),
    .A2(_02814_),
    .A3(_02825_),
    .B1(_01452_),
    .X(_02859_));
 sky130_fd_sc_hd__o221a_2 _07939_ (.A1(_01065_),
    .A2(_01074_),
    .B1(_01870_),
    .B2(_02849_),
    .C1(_02798_),
    .X(_02860_));
 sky130_fd_sc_hd__o22ai_2 _07940_ (.A1(_02858_),
    .A2(_02859_),
    .B1(_02803_),
    .B2(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__o2111a_2 _07941_ (.A1(_02851_),
    .A2(_02803_),
    .B1(_02856_),
    .C1(_02751_),
    .D1(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__nor2_2 _07942_ (.A(\rvsingle.dp.rf.rf[0][0] ),
    .B(_01256_),
    .Y(_02863_));
 sky130_fd_sc_hd__and2b_2 _07943_ (.A_N(\rvsingle.dp.rf.rf[1][0] ),
    .B(_01675_),
    .X(_02864_));
 sky130_fd_sc_hd__o21a_2 _07944_ (.A1(\rvsingle.dp.rf.rf[2][0] ),
    .A2(_01753_),
    .B1(_01596_),
    .X(_02865_));
 sky130_fd_sc_hd__o21ai_2 _07945_ (.A1(\rvsingle.dp.rf.rf[3][0] ),
    .A2(_01842_),
    .B1(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__o311a_2 _07946_ (.A1(_01648_),
    .A2(_02863_),
    .A3(_02864_),
    .B1(_01600_),
    .C1(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__nor2_2 _07947_ (.A(\rvsingle.dp.rf.rf[4][0] ),
    .B(_01643_),
    .Y(_02868_));
 sky130_fd_sc_hd__o21ai_2 _07948_ (.A1(\rvsingle.dp.rf.rf[5][0] ),
    .A2(_01796_),
    .B1(_01092_),
    .Y(_02869_));
 sky130_fd_sc_hd__o21a_2 _07949_ (.A1(\rvsingle.dp.rf.rf[6][0] ),
    .A2(_01675_),
    .B1(_01596_),
    .X(_02870_));
 sky130_fd_sc_hd__o21ai_2 _07950_ (.A1(\rvsingle.dp.rf.rf[7][0] ),
    .A2(_01842_),
    .B1(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__o211a_2 _07951_ (.A1(_02868_),
    .A2(_02869_),
    .B1(_01617_),
    .C1(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__inv_2 _07952_ (.A(net248),
    .Y(_02873_));
 sky130_fd_sc_hd__o21ai_2 _07953_ (.A1(\rvsingle.dp.rf.rf[10][0] ),
    .A2(_01493_),
    .B1(_01552_),
    .Y(_02874_));
 sky130_fd_sc_hd__a21oi_2 _07954_ (.A1(_02873_),
    .A2(_01848_),
    .B1(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__inv_2 _07955_ (.A(\rvsingle.dp.rf.rf[9][0] ),
    .Y(_02876_));
 sky130_fd_sc_hd__nor2_2 _07956_ (.A(\rvsingle.dp.rf.rf[8][0] ),
    .B(_01619_),
    .Y(_02877_));
 sky130_fd_sc_hd__a211oi_2 _07957_ (.A1(_02876_),
    .A2(_01643_),
    .B1(_01105_),
    .C1(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__nor2_2 _07958_ (.A(\rvsingle.dp.rf.rf[14][0] ),
    .B(_01518_),
    .Y(_02879_));
 sky130_fd_sc_hd__o21ai_2 _07959_ (.A1(\rvsingle.dp.rf.rf[15][0] ),
    .A2(_02478_),
    .B1(_01490_),
    .Y(_02880_));
 sky130_fd_sc_hd__nor2_2 _07960_ (.A(\rvsingle.dp.rf.rf[12][0] ),
    .B(_01619_),
    .Y(_02881_));
 sky130_fd_sc_hd__o21ai_2 _07961_ (.A1(\rvsingle.dp.rf.rf[13][0] ),
    .A2(_01487_),
    .B1(_01496_),
    .Y(_02882_));
 sky130_fd_sc_hd__o221ai_2 _07962_ (.A1(_02879_),
    .A2(_02880_),
    .B1(_02881_),
    .B2(_02882_),
    .C1(_02488_),
    .Y(_02883_));
 sky130_fd_sc_hd__o311ai_2 _07963_ (.A1(_01503_),
    .A2(_02875_),
    .A3(_02878_),
    .B1(_01116_),
    .C1(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__o311ai_2 _07964_ (.A1(_01526_),
    .A2(_02867_),
    .A3(_02872_),
    .B1(_02884_),
    .C1(_01593_),
    .Y(_02885_));
 sky130_fd_sc_hd__nor2_2 _07965_ (.A(\rvsingle.dp.rf.rf[28][0] ),
    .B(_01126_),
    .Y(_02886_));
 sky130_fd_sc_hd__o21ai_2 _07966_ (.A1(\rvsingle.dp.rf.rf[29][0] ),
    .A2(_01796_),
    .B1(_02485_),
    .Y(_02887_));
 sky130_fd_sc_hd__o21a_2 _07967_ (.A1(\rvsingle.dp.rf.rf[30][0] ),
    .A2(_01642_),
    .B1(_01596_),
    .X(_02888_));
 sky130_fd_sc_hd__o21ai_2 _07968_ (.A1(\rvsingle.dp.rf.rf[31][0] ),
    .A2(_01646_),
    .B1(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__o211a_2 _07969_ (.A1(_02886_),
    .A2(_02887_),
    .B1(_01617_),
    .C1(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__o21ba_2 _07970_ (.A1(\rvsingle.dp.rf.rf[24][0] ),
    .A2(_02005_),
    .B1_N(_01530_),
    .X(_02891_));
 sky130_fd_sc_hd__o21ai_2 _07971_ (.A1(\rvsingle.dp.rf.rf[25][0] ),
    .A2(_01796_),
    .B1(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__or2b_2 _07972_ (.A(\rvsingle.dp.rf.rf[27][0] ),
    .B_N(_01561_),
    .X(_02893_));
 sky130_fd_sc_hd__o211ai_2 _07973_ (.A1(\rvsingle.dp.rf.rf[26][0] ),
    .A2(_01562_),
    .B1(_02320_),
    .C1(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__a31o_2 _07974_ (.A1(_01600_),
    .A2(_02892_),
    .A3(_02894_),
    .B1(_02364_),
    .X(_02895_));
 sky130_fd_sc_hd__nor2_2 _07975_ (.A(\rvsingle.dp.rf.rf[16][0] ),
    .B(_01603_),
    .Y(_02896_));
 sky130_fd_sc_hd__o21ai_2 _07976_ (.A1(\rvsingle.dp.rf.rf[17][0] ),
    .A2(_01677_),
    .B1(_02485_),
    .Y(_02897_));
 sky130_fd_sc_hd__nor2_2 _07977_ (.A(\rvsingle.dp.rf.rf[18][0] ),
    .B(_01126_),
    .Y(_02898_));
 sky130_fd_sc_hd__o21ai_2 _07978_ (.A1(\rvsingle.dp.rf.rf[19][0] ),
    .A2(_01677_),
    .B1(_01531_),
    .Y(_02899_));
 sky130_fd_sc_hd__o221a_2 _07979_ (.A1(_02896_),
    .A2(_02897_),
    .B1(_02898_),
    .B2(_02899_),
    .C1(_01600_),
    .X(_02900_));
 sky130_fd_sc_hd__or2_2 _07980_ (.A(\rvsingle.dp.rf.rf[20][0] ),
    .B(_01255_),
    .X(_02901_));
 sky130_fd_sc_hd__o211ai_2 _07981_ (.A1(\rvsingle.dp.rf.rf[21][0] ),
    .A2(_01796_),
    .B1(_02485_),
    .C1(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__o21a_2 _07982_ (.A1(\rvsingle.dp.rf.rf[22][0] ),
    .A2(_01797_),
    .B1(_01104_),
    .X(_02903_));
 sky130_fd_sc_hd__o21ai_2 _07983_ (.A1(\rvsingle.dp.rf.rf[23][0] ),
    .A2(_01646_),
    .B1(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__a31o_2 _07984_ (.A1(_02902_),
    .A2(_01617_),
    .A3(_02904_),
    .B1(_02491_),
    .X(_02905_));
 sky130_fd_sc_hd__o221ai_2 _07985_ (.A1(_02890_),
    .A2(_02895_),
    .B1(_02900_),
    .B2(_02905_),
    .C1(_01682_),
    .Y(_02906_));
 sky130_fd_sc_hd__a31oi_2 _07986_ (.A1(_01592_),
    .A2(_02885_),
    .A3(_02906_),
    .B1(_01178_),
    .Y(_02907_));
 sky130_fd_sc_hd__buf_1 _07987_ (.A(_01081_),
    .X(_02908_));
 sky130_fd_sc_hd__buf_1 _07988_ (.A(Instr[3]),
    .X(_02909_));
 sky130_fd_sc_hd__buf_1 _07989_ (.A(Instr[2]),
    .X(_02910_));
 sky130_fd_sc_hd__nor4_2 _07990_ (.A(_01067_),
    .B(_02909_),
    .C(_02910_),
    .D(_01173_),
    .Y(_02911_));
 sky130_fd_sc_hd__buf_1 _07991_ (.A(_01076_),
    .X(_02912_));
 sky130_fd_sc_hd__o211ai_2 _07992_ (.A1(_01175_),
    .A2(_02911_),
    .B1(Instr[7]),
    .C1(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__o211ai_2 _07993_ (.A1(_01067_),
    .A2(_01078_),
    .B1(_01080_),
    .C1(_01099_),
    .Y(_02914_));
 sky130_fd_sc_hd__a22oi_2 _07994_ (.A1(_02908_),
    .A2(_01067_),
    .B1(_02913_),
    .B2(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__nor2_2 _07995_ (.A(_01903_),
    .B(\rvsingle.dp.rf.rf[26][0] ),
    .Y(_02916_));
 sky130_fd_sc_hd__and2b_2 _07996_ (.A_N(\rvsingle.dp.rf.rf[27][0] ),
    .B(_01240_),
    .X(_02917_));
 sky130_fd_sc_hd__o21ba_2 _07997_ (.A1(_01425_),
    .A2(\rvsingle.dp.rf.rf[24][0] ),
    .B1_N(_01197_),
    .X(_02918_));
 sky130_fd_sc_hd__o21ai_2 _07998_ (.A1(_01423_),
    .A2(\rvsingle.dp.rf.rf[25][0] ),
    .B1(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__o31ai_2 _07999_ (.A1(_01307_),
    .A2(_02916_),
    .A3(_02917_),
    .B1(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__nor2_2 _08000_ (.A(_01416_),
    .B(\rvsingle.dp.rf.rf[30][0] ),
    .Y(_02921_));
 sky130_fd_sc_hd__o21ai_2 _08001_ (.A1(\rvsingle.dp.rf.rf[31][0] ),
    .A2(_01423_),
    .B1(_01427_),
    .Y(_02922_));
 sky130_fd_sc_hd__or2_2 _08002_ (.A(_01327_),
    .B(\rvsingle.dp.rf.rf[28][0] ),
    .X(_02923_));
 sky130_fd_sc_hd__o211ai_2 _08003_ (.A1(\rvsingle.dp.rf.rf[29][0] ),
    .A2(_01423_),
    .B1(_01307_),
    .C1(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__o211ai_2 _08004_ (.A1(_02921_),
    .A2(_02922_),
    .B1(_01172_),
    .C1(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__o211ai_2 _08005_ (.A1(_02273_),
    .A2(_02920_),
    .B1(_02925_),
    .C1(_01446_),
    .Y(_02926_));
 sky130_fd_sc_hd__nor2_2 _08006_ (.A(_02450_),
    .B(\rvsingle.dp.rf.rf[16][0] ),
    .Y(_02927_));
 sky130_fd_sc_hd__o21bai_2 _08007_ (.A1(\rvsingle.dp.rf.rf[17][0] ),
    .A2(_01423_),
    .B1_N(_01454_),
    .Y(_02928_));
 sky130_fd_sc_hd__buf_1 _08008_ (.A(_01293_),
    .X(_02929_));
 sky130_fd_sc_hd__o21a_2 _08009_ (.A1(_01240_),
    .A2(\rvsingle.dp.rf.rf[18][0] ),
    .B1(_01197_),
    .X(_02930_));
 sky130_fd_sc_hd__o21ai_2 _08010_ (.A1(\rvsingle.dp.rf.rf[19][0] ),
    .A2(_02929_),
    .B1(_02930_),
    .Y(_02931_));
 sky130_fd_sc_hd__o211ai_2 _08011_ (.A1(_02927_),
    .A2(_02928_),
    .B1(_01206_),
    .C1(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__or2_2 _08012_ (.A(_01327_),
    .B(\rvsingle.dp.rf.rf[20][0] ),
    .X(_02933_));
 sky130_fd_sc_hd__o211ai_2 _08013_ (.A1(\rvsingle.dp.rf.rf[21][0] ),
    .A2(_02929_),
    .B1(_01307_),
    .C1(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__o21a_2 _08014_ (.A1(_01425_),
    .A2(\rvsingle.dp.rf.rf[22][0] ),
    .B1(_01197_),
    .X(_02935_));
 sky130_fd_sc_hd__o21ai_2 _08015_ (.A1(\rvsingle.dp.rf.rf[23][0] ),
    .A2(_02929_),
    .B1(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand3_2 _08016_ (.A(_02934_),
    .B(_01172_),
    .C(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand3_2 _08017_ (.A(_01217_),
    .B(_02932_),
    .C(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__nand3_2 _08018_ (.A(_02926_),
    .B(_02938_),
    .C(_01187_),
    .Y(_02939_));
 sky130_fd_sc_hd__o21bai_2 _08019_ (.A1(_01725_),
    .A2(\rvsingle.dp.rf.rf[8][0] ),
    .B1_N(_01454_),
    .Y(_02940_));
 sky130_fd_sc_hd__a21oi_2 _08020_ (.A1(_02876_),
    .A2(_01691_),
    .B1(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__o21ai_2 _08021_ (.A1(_02440_),
    .A2(\rvsingle.dp.rf.rf[10][0] ),
    .B1(_01243_),
    .Y(_02942_));
 sky130_fd_sc_hd__a21oi_2 _08022_ (.A1(_02873_),
    .A2(_01707_),
    .B1(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__nor2_2 _08023_ (.A(_01328_),
    .B(\rvsingle.dp.rf.rf[14][0] ),
    .Y(_02944_));
 sky130_fd_sc_hd__o21ai_2 _08024_ (.A1(\rvsingle.dp.rf.rf[15][0] ),
    .A2(_01294_),
    .B1(_01243_),
    .Y(_02945_));
 sky130_fd_sc_hd__or2_2 _08025_ (.A(_01327_),
    .B(\rvsingle.dp.rf.rf[12][0] ),
    .X(_02946_));
 sky130_fd_sc_hd__o211ai_2 _08026_ (.A1(\rvsingle.dp.rf.rf[13][0] ),
    .A2(_01423_),
    .B1(_01307_),
    .C1(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__o211ai_2 _08027_ (.A1(_02944_),
    .A2(_02945_),
    .B1(_01172_),
    .C1(_02947_),
    .Y(_02948_));
 sky130_fd_sc_hd__o311ai_2 _08028_ (.A1(_01444_),
    .A2(_02941_),
    .A3(_02943_),
    .B1(_01215_),
    .C1(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__o21bai_2 _08029_ (.A1(\rvsingle.dp.rf.rf[0][0] ),
    .A2(_02440_),
    .B1_N(_01454_),
    .Y(_02950_));
 sky130_fd_sc_hd__and2b_2 _08030_ (.A_N(\rvsingle.dp.rf.rf[1][0] ),
    .B(_01690_),
    .X(_02951_));
 sky130_fd_sc_hd__o21ai_2 _08031_ (.A1(_02950_),
    .A2(_02951_),
    .B1(_01206_),
    .Y(_02952_));
 sky130_fd_sc_hd__or2_2 _08032_ (.A(_01425_),
    .B(\rvsingle.dp.rf.rf[2][0] ),
    .X(_02953_));
 sky130_fd_sc_hd__o211a_2 _08033_ (.A1(_01423_),
    .A2(\rvsingle.dp.rf.rf[3][0] ),
    .B1(_01427_),
    .C1(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__nor2_2 _08034_ (.A(_02176_),
    .B(\rvsingle.dp.rf.rf[4][0] ),
    .Y(_02955_));
 sky130_fd_sc_hd__o21ai_2 _08035_ (.A1(\rvsingle.dp.rf.rf[5][0] ),
    .A2(_01423_),
    .B1(_01307_),
    .Y(_02956_));
 sky130_fd_sc_hd__o21a_2 _08036_ (.A1(_01240_),
    .A2(\rvsingle.dp.rf.rf[6][0] ),
    .B1(_01454_),
    .X(_02957_));
 sky130_fd_sc_hd__o21ai_2 _08037_ (.A1(\rvsingle.dp.rf.rf[7][0] ),
    .A2(_02929_),
    .B1(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__o211ai_2 _08038_ (.A1(_02955_),
    .A2(_02956_),
    .B1(_01172_),
    .C1(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__o211ai_2 _08039_ (.A1(_02952_),
    .A2(_02954_),
    .B1(_01216_),
    .C1(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__nand3_2 _08040_ (.A(_01315_),
    .B(_02949_),
    .C(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__o311a_2 _08041_ (.A1(_01337_),
    .A2(_01451_),
    .A3(_01245_),
    .B1(_02939_),
    .C1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__o21ai_2 _08042_ (.A1(_01870_),
    .A2(_02915_),
    .B1(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__nand4_2 _08043_ (.A(_02885_),
    .B(_01481_),
    .C(_01592_),
    .D(_02906_),
    .Y(_02964_));
 sky130_fd_sc_hd__a221o_2 _08044_ (.A1(_01067_),
    .A2(_01081_),
    .B1(_02914_),
    .B2(_02913_),
    .C1(_01083_),
    .X(_02965_));
 sky130_fd_sc_hd__nand3_2 _08045_ (.A(_02964_),
    .B(_02965_),
    .C(_01183_),
    .Y(_02966_));
 sky130_fd_sc_hd__o21ai_2 _08046_ (.A1(_02907_),
    .A2(_02963_),
    .B1(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__or2_2 _08047_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[10][1] ),
    .X(_02968_));
 sky130_fd_sc_hd__o211a_2 _08048_ (.A1(_01440_),
    .A2(\rvsingle.dp.rf.rf[11][1] ),
    .B1(_02162_),
    .C1(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__or2_2 _08049_ (.A(_01690_),
    .B(\rvsingle.dp.rf.rf[8][1] ),
    .X(_02970_));
 sky130_fd_sc_hd__o211ai_2 _08050_ (.A1(\rvsingle.dp.rf.rf[9][1] ),
    .A2(_02271_),
    .B1(_02268_),
    .C1(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__nand2_2 _08051_ (.A(_01460_),
    .B(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__mux4_2 _08052_ (.A0(\rvsingle.dp.rf.rf[12][1] ),
    .A1(\rvsingle.dp.rf.rf[13][1] ),
    .A2(\rvsingle.dp.rf.rf[14][1] ),
    .A3(\rvsingle.dp.rf.rf[15][1] ),
    .S0(_01903_),
    .S1(_01470_),
    .X(_02973_));
 sky130_fd_sc_hd__o221ai_2 _08053_ (.A1(_02969_),
    .A2(_02972_),
    .B1(_01207_),
    .B2(_02973_),
    .C1(_02438_),
    .Y(_02974_));
 sky130_fd_sc_hd__mux4_2 _08054_ (.A0(\rvsingle.dp.rf.rf[0][1] ),
    .A1(\rvsingle.dp.rf.rf[1][1] ),
    .A2(\rvsingle.dp.rf.rf[2][1] ),
    .A3(\rvsingle.dp.rf.rf[3][1] ),
    .S0(_02440_),
    .S1(_01470_),
    .X(_02975_));
 sky130_fd_sc_hd__nor2_2 _08055_ (.A(_01695_),
    .B(\rvsingle.dp.rf.rf[4][1] ),
    .Y(_02976_));
 sky130_fd_sc_hd__o21ai_2 _08056_ (.A1(\rvsingle.dp.rf.rf[5][1] ),
    .A2(_02271_),
    .B1(_01436_),
    .Y(_02977_));
 sky130_fd_sc_hd__o21a_2 _08057_ (.A1(_01468_),
    .A2(\rvsingle.dp.rf.rf[6][1] ),
    .B1(_01198_),
    .X(_02978_));
 sky130_fd_sc_hd__o21ai_2 _08058_ (.A1(\rvsingle.dp.rf.rf[7][1] ),
    .A2(_01295_),
    .B1(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__o211ai_2 _08059_ (.A1(_02976_),
    .A2(_02977_),
    .B1(_02273_),
    .C1(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__o211ai_2 _08060_ (.A1(_01229_),
    .A2(_02975_),
    .B1(_02980_),
    .C1(_02447_),
    .Y(_02981_));
 sky130_fd_sc_hd__nand2_2 _08061_ (.A(_02974_),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__mux2_2 _08062_ (.A0(\rvsingle.dp.rf.rf[16][1] ),
    .A1(\rvsingle.dp.rf.rf[17][1] ),
    .S(_01241_),
    .X(_02983_));
 sky130_fd_sc_hd__or2_2 _08063_ (.A(_01191_),
    .B(\rvsingle.dp.rf.rf[18][1] ),
    .X(_02984_));
 sky130_fd_sc_hd__o211a_2 _08064_ (.A1(_02275_),
    .A2(\rvsingle.dp.rf.rf[19][1] ),
    .B1(_02162_),
    .C1(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__a211oi_2 _08065_ (.A1(_02983_),
    .A2(_01437_),
    .B1(_01702_),
    .C1(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__mux4_2 _08066_ (.A0(\rvsingle.dp.rf.rf[20][1] ),
    .A1(\rvsingle.dp.rf.rf[21][1] ),
    .A2(\rvsingle.dp.rf.rf[22][1] ),
    .A3(\rvsingle.dp.rf.rf[23][1] ),
    .S0(_02440_),
    .S1(_01470_),
    .X(_02987_));
 sky130_fd_sc_hd__o21ai_2 _08067_ (.A1(_01207_),
    .A2(_02987_),
    .B1(_02447_),
    .Y(_02988_));
 sky130_fd_sc_hd__mux4_2 _08068_ (.A0(\rvsingle.dp.rf.rf[24][1] ),
    .A1(\rvsingle.dp.rf.rf[25][1] ),
    .A2(\rvsingle.dp.rf.rf[26][1] ),
    .A3(\rvsingle.dp.rf.rf[27][1] ),
    .S0(_01903_),
    .S1(_01470_),
    .X(_02989_));
 sky130_fd_sc_hd__nor2_2 _08069_ (.A(_01695_),
    .B(\rvsingle.dp.rf.rf[30][1] ),
    .Y(_02990_));
 sky130_fd_sc_hd__o21ai_2 _08070_ (.A1(\rvsingle.dp.rf.rf[31][1] ),
    .A2(_01440_),
    .B1(_02162_),
    .Y(_02991_));
 sky130_fd_sc_hd__or2_2 _08071_ (.A(_01349_),
    .B(\rvsingle.dp.rf.rf[28][1] ),
    .X(_02992_));
 sky130_fd_sc_hd__o211ai_2 _08072_ (.A1(\rvsingle.dp.rf.rf[29][1] ),
    .A2(_02275_),
    .B1(_01436_),
    .C1(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__o211ai_2 _08073_ (.A1(_02990_),
    .A2(_02991_),
    .B1(_02273_),
    .C1(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__o211ai_2 _08074_ (.A1(_02302_),
    .A2(_02989_),
    .B1(_02994_),
    .C1(_02438_),
    .Y(_02995_));
 sky130_fd_sc_hd__o211ai_2 _08075_ (.A1(_02986_),
    .A2(_02988_),
    .B1(_01187_),
    .C1(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hd__o21ai_2 _08076_ (.A1(_01188_),
    .A2(_02982_),
    .B1(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__nor2_2 _08077_ (.A(_01847_),
    .B(\rvsingle.dp.rf.rf[2][1] ),
    .Y(_02998_));
 sky130_fd_sc_hd__o21ai_2 _08078_ (.A1(\rvsingle.dp.rf.rf[3][1] ),
    .A2(_01645_),
    .B1(_01596_),
    .Y(_02999_));
 sky130_fd_sc_hd__or2b_2 _08079_ (.A(\rvsingle.dp.rf.rf[1][1] ),
    .B_N(_01124_),
    .X(_03000_));
 sky130_fd_sc_hd__o211ai_2 _08080_ (.A1(_01797_),
    .A2(\rvsingle.dp.rf.rf[0][1] ),
    .B1(_03000_),
    .C1(_01667_),
    .Y(_03001_));
 sky130_fd_sc_hd__o211a_2 _08081_ (.A1(_02998_),
    .A2(_02999_),
    .B1(_03001_),
    .C1(_01564_),
    .X(_03002_));
 sky130_fd_sc_hd__or2b_2 _08082_ (.A(\rvsingle.dp.rf.rf[5][1] ),
    .B_N(_01606_),
    .X(_03003_));
 sky130_fd_sc_hd__o211ai_2 _08083_ (.A1(_01642_),
    .A2(\rvsingle.dp.rf.rf[4][1] ),
    .B1(_03003_),
    .C1(_01667_),
    .Y(_03004_));
 sky130_fd_sc_hd__or2b_2 _08084_ (.A(\rvsingle.dp.rf.rf[7][1] ),
    .B_N(_01606_),
    .X(_03005_));
 sky130_fd_sc_hd__o211ai_2 _08085_ (.A1(_01797_),
    .A2(\rvsingle.dp.rf.rf[6][1] ),
    .B1(_01647_),
    .C1(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__a31o_2 _08086_ (.A1(_03004_),
    .A2(_03006_),
    .A3(_01502_),
    .B1(_01115_),
    .X(_03007_));
 sky130_fd_sc_hd__nor2_2 _08087_ (.A(_01797_),
    .B(\rvsingle.dp.rf.rf[10][1] ),
    .Y(_03008_));
 sky130_fd_sc_hd__o21ai_2 _08088_ (.A1(\rvsingle.dp.rf.rf[11][1] ),
    .A2(_01645_),
    .B1(_01647_),
    .Y(_03009_));
 sky130_fd_sc_hd__nor2_2 _08089_ (.A(_01642_),
    .B(\rvsingle.dp.rf.rf[8][1] ),
    .Y(_03010_));
 sky130_fd_sc_hd__o21ai_2 _08090_ (.A1(\rvsingle.dp.rf.rf[9][1] ),
    .A2(_01645_),
    .B1(_01667_),
    .Y(_03011_));
 sky130_fd_sc_hd__o221ai_2 _08091_ (.A1(_03008_),
    .A2(_03009_),
    .B1(_03010_),
    .B2(_03011_),
    .C1(_01564_),
    .Y(_03012_));
 sky130_fd_sc_hd__or2_2 _08092_ (.A(_01606_),
    .B(\rvsingle.dp.rf.rf[12][1] ),
    .X(_03013_));
 sky130_fd_sc_hd__o211ai_2 _08093_ (.A1(\rvsingle.dp.rf.rf[13][1] ),
    .A2(_01087_),
    .B1(_01667_),
    .C1(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__o21a_2 _08094_ (.A1(_01096_),
    .A2(\rvsingle.dp.rf.rf[14][1] ),
    .B1(_01610_),
    .X(_03015_));
 sky130_fd_sc_hd__o21ai_2 _08095_ (.A1(\rvsingle.dp.rf.rf[15][1] ),
    .A2(_01087_),
    .B1(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__nand3_2 _08096_ (.A(_03014_),
    .B(_01502_),
    .C(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__nand3_2 _08097_ (.A(_03012_),
    .B(_02491_),
    .C(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__o211ai_2 _08098_ (.A1(_03002_),
    .A2(_03007_),
    .B1(_01376_),
    .C1(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__nor2_2 _08099_ (.A(_01602_),
    .B(\rvsingle.dp.rf.rf[20][1] ),
    .Y(_03020_));
 sky130_fd_sc_hd__and2b_2 _08100_ (.A_N(\rvsingle.dp.rf.rf[21][1] ),
    .B(_01381_),
    .X(_03021_));
 sky130_fd_sc_hd__or2b_2 _08101_ (.A(\rvsingle.dp.rf.rf[23][1] ),
    .B_N(_01124_),
    .X(_03022_));
 sky130_fd_sc_hd__o211ai_2 _08102_ (.A1(_01769_),
    .A2(\rvsingle.dp.rf.rf[22][1] ),
    .B1(_01604_),
    .C1(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__o311ai_2 _08103_ (.A1(_01880_),
    .A2(_03020_),
    .A3(_03021_),
    .B1(_01110_),
    .C1(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__nor2_2 _08104_ (.A(_01602_),
    .B(\rvsingle.dp.rf.rf[16][1] ),
    .Y(_03025_));
 sky130_fd_sc_hd__and2b_2 _08105_ (.A_N(\rvsingle.dp.rf.rf[17][1] ),
    .B(_01381_),
    .X(_03026_));
 sky130_fd_sc_hd__or2b_2 _08106_ (.A(\rvsingle.dp.rf.rf[19][1] ),
    .B_N(_01124_),
    .X(_03027_));
 sky130_fd_sc_hd__o211ai_2 _08107_ (.A1(_01769_),
    .A2(\rvsingle.dp.rf.rf[18][1] ),
    .B1(_01604_),
    .C1(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__o311ai_2 _08108_ (.A1(_01880_),
    .A2(_03025_),
    .A3(_03026_),
    .B1(_01599_),
    .C1(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__nand3_2 _08109_ (.A(_02364_),
    .B(_03024_),
    .C(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__nor2_2 _08110_ (.A(_01602_),
    .B(\rvsingle.dp.rf.rf[24][1] ),
    .Y(_03031_));
 sky130_fd_sc_hd__and2b_2 _08111_ (.A_N(\rvsingle.dp.rf.rf[25][1] ),
    .B(_01381_),
    .X(_03032_));
 sky130_fd_sc_hd__or2b_2 _08112_ (.A(\rvsingle.dp.rf.rf[27][1] ),
    .B_N(_01124_),
    .X(_03033_));
 sky130_fd_sc_hd__o211ai_2 _08113_ (.A1(_01650_),
    .A2(\rvsingle.dp.rf.rf[26][1] ),
    .B1(_01104_),
    .C1(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__o311ai_2 _08114_ (.A1(_01259_),
    .A2(_03031_),
    .A3(_03032_),
    .B1(_01599_),
    .C1(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__and2b_2 _08115_ (.A_N(\rvsingle.dp.rf.rf[29][1] ),
    .B(_01544_),
    .X(_03036_));
 sky130_fd_sc_hd__o21ai_2 _08116_ (.A1(_01769_),
    .A2(\rvsingle.dp.rf.rf[28][1] ),
    .B1(_01091_),
    .Y(_03037_));
 sky130_fd_sc_hd__or2b_2 _08117_ (.A(\rvsingle.dp.rf.rf[31][1] ),
    .B_N(_01124_),
    .X(_03038_));
 sky130_fd_sc_hd__o211ai_2 _08118_ (.A1(_02005_),
    .A2(\rvsingle.dp.rf.rf[30][1] ),
    .B1(_01104_),
    .C1(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__o211ai_2 _08119_ (.A1(_03036_),
    .A2(_03037_),
    .B1(_01502_),
    .C1(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__nand3_2 _08120_ (.A(_03035_),
    .B(_01115_),
    .C(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__nand3_2 _08121_ (.A(_03030_),
    .B(_01145_),
    .C(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__nand4_2 _08122_ (.A(_03019_),
    .B(_01082_),
    .C(_01152_),
    .D(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand4_2 _08123_ (.A(Instr[8]),
    .B(_01076_),
    .C(_01071_),
    .D(_01062_),
    .Y(_03044_));
 sky130_fd_sc_hd__o21ai_2 _08124_ (.A1(_01856_),
    .A2(_01069_),
    .B1(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand2_2 _08125_ (.A(_01177_),
    .B(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__a21oi_2 _08126_ (.A1(_03043_),
    .A2(_03046_),
    .B1(_01485_),
    .Y(_03047_));
 sky130_fd_sc_hd__o211a_2 _08127_ (.A1(_01065_),
    .A2(_01074_),
    .B1(_03043_),
    .C1(_03046_),
    .X(_03048_));
 sky130_fd_sc_hd__o22ai_2 _08128_ (.A1(_01452_),
    .A2(_02997_),
    .B1(_03047_),
    .B2(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__o211a_2 _08129_ (.A1(_02315_),
    .A2(_02982_),
    .B1(_02996_),
    .C1(_01246_),
    .X(_03050_));
 sky130_fd_sc_hd__o211ai_2 _08130_ (.A1(_02473_),
    .A2(_02318_),
    .B1(_03043_),
    .C1(_03046_),
    .Y(_03051_));
 sky130_fd_sc_hd__nand2_2 _08131_ (.A(_03050_),
    .B(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__o2bb2ai_2 _08132_ (.A1_N(_02967_),
    .A2_N(_03049_),
    .B1(_03047_),
    .B2(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__a22oi_2 _08133_ (.A1(_02751_),
    .A2(_02857_),
    .B1(_02862_),
    .B2(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__a21o_2 _08134_ (.A1(_02530_),
    .A2(_02533_),
    .B1(_01591_),
    .X(_03055_));
 sky130_fd_sc_hd__nand3_2 _08135_ (.A(_03055_),
    .B(_02572_),
    .C(_02570_),
    .Y(_03056_));
 sky130_fd_sc_hd__a2bb2oi_2 _08136_ (.A1_N(_02469_),
    .A2_N(_02608_),
    .B1(_02666_),
    .B2(_02664_),
    .Y(_03057_));
 sky130_fd_sc_hd__a21oi_2 _08137_ (.A1(_03056_),
    .A2(_02667_),
    .B1(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__a31o_2 _08138_ (.A1(_01592_),
    .A2(_02346_),
    .A3(_02371_),
    .B1(_01178_),
    .X(_03059_));
 sky130_fd_sc_hd__o211ai_2 _08139_ (.A1(Instr[27]),
    .A2(_01084_),
    .B1(_01584_),
    .C1(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__a21oi_2 _08140_ (.A1(_03060_),
    .A2(_02373_),
    .B1(_02317_),
    .Y(_03061_));
 sky130_fd_sc_hd__o22ai_2 _08141_ (.A1(_02377_),
    .A2(_02374_),
    .B1(_02464_),
    .B2(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__a21oi_2 _08142_ (.A1(_02476_),
    .A2(_03058_),
    .B1(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__o21ai_2 _08143_ (.A1(_02668_),
    .A2(_03054_),
    .B1(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__nor2_2 _08144_ (.A(_01382_),
    .B(\rvsingle.dp.rf.rf[18][11] ),
    .Y(_03065_));
 sky130_fd_sc_hd__o21ai_2 _08145_ (.A1(\rvsingle.dp.rf.rf[19][11] ),
    .A2(_01860_),
    .B1(_01259_),
    .Y(_03066_));
 sky130_fd_sc_hd__o21ba_2 _08146_ (.A1(_01779_),
    .A2(\rvsingle.dp.rf.rf[16][11] ),
    .B1_N(_01610_),
    .X(_03067_));
 sky130_fd_sc_hd__o21ai_2 _08147_ (.A1(_02379_),
    .A2(\rvsingle.dp.rf.rf[17][11] ),
    .B1(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__o211ai_2 _08148_ (.A1(_03065_),
    .A2(_03066_),
    .B1(_03068_),
    .C1(_01131_),
    .Y(_03069_));
 sky130_fd_sc_hd__nor2_2 _08149_ (.A(_01382_),
    .B(\rvsingle.dp.rf.rf[20][11] ),
    .Y(_03070_));
 sky130_fd_sc_hd__o21bai_2 _08150_ (.A1(\rvsingle.dp.rf.rf[21][11] ),
    .A2(_01860_),
    .B1_N(_01530_),
    .Y(_03071_));
 sky130_fd_sc_hd__o21a_2 _08151_ (.A1(_01498_),
    .A2(\rvsingle.dp.rf.rf[22][11] ),
    .B1(_01519_),
    .X(_03072_));
 sky130_fd_sc_hd__o21ai_2 _08152_ (.A1(\rvsingle.dp.rf.rf[23][11] ),
    .A2(_01539_),
    .B1(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__o211ai_2 _08153_ (.A1(_03070_),
    .A2(_03071_),
    .B1(_02323_),
    .C1(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand3_2 _08154_ (.A(_01156_),
    .B(_03069_),
    .C(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__o21bai_2 _08155_ (.A1(_01743_),
    .A2(\rvsingle.dp.rf.rf[24][11] ),
    .B1_N(_01519_),
    .Y(_03076_));
 sky130_fd_sc_hd__and2b_2 _08156_ (.A_N(\rvsingle.dp.rf.rf[25][11] ),
    .B(_01492_),
    .X(_03077_));
 sky130_fd_sc_hd__o21ai_2 _08157_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_01564_),
    .Y(_03078_));
 sky130_fd_sc_hd__or2b_2 _08158_ (.A(\rvsingle.dp.rf.rf[27][11] ),
    .B_N(_01566_),
    .X(_03079_));
 sky130_fd_sc_hd__o211a_2 _08159_ (.A1(_01630_),
    .A2(\rvsingle.dp.rf.rf[26][11] ),
    .B1(_01259_),
    .C1(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__o21ba_2 _08160_ (.A1(_01779_),
    .A2(\rvsingle.dp.rf.rf[28][11] ),
    .B1_N(_01610_),
    .X(_03081_));
 sky130_fd_sc_hd__o21ai_2 _08161_ (.A1(_02379_),
    .A2(\rvsingle.dp.rf.rf[29][11] ),
    .B1(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__o21a_2 _08162_ (.A1(_01544_),
    .A2(\rvsingle.dp.rf.rf[30][11] ),
    .B1(_01258_),
    .X(_03083_));
 sky130_fd_sc_hd__o21ai_2 _08163_ (.A1(\rvsingle.dp.rf.rf[31][11] ),
    .A2(_01860_),
    .B1(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__nand3_2 _08164_ (.A(_03082_),
    .B(_01111_),
    .C(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__o211ai_2 _08165_ (.A1(_03078_),
    .A2(_03080_),
    .B1(_03085_),
    .C1(_02491_),
    .Y(_03086_));
 sky130_fd_sc_hd__nand3_2 _08166_ (.A(_03075_),
    .B(_01146_),
    .C(_03086_),
    .Y(_03087_));
 sky130_fd_sc_hd__nor2_2 _08167_ (.A(_01097_),
    .B(\rvsingle.dp.rf.rf[4][11] ),
    .Y(_03088_));
 sky130_fd_sc_hd__and2b_2 _08168_ (.A_N(\rvsingle.dp.rf.rf[5][11] ),
    .B(_01613_),
    .X(_03089_));
 sky130_fd_sc_hd__or2_2 _08169_ (.A(_01381_),
    .B(\rvsingle.dp.rf.rf[6][11] ),
    .X(_03090_));
 sky130_fd_sc_hd__o211ai_2 _08170_ (.A1(_02379_),
    .A2(\rvsingle.dp.rf.rf[7][11] ),
    .B1(_02031_),
    .C1(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__o311a_2 _08171_ (.A1(_01552_),
    .A2(_03088_),
    .A3(_03089_),
    .B1(_02323_),
    .C1(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__o21bai_2 _08172_ (.A1(_02005_),
    .A2(\rvsingle.dp.rf.rf[0][11] ),
    .B1_N(_01519_),
    .Y(_03093_));
 sky130_fd_sc_hd__and2b_2 _08173_ (.A_N(\rvsingle.dp.rf.rf[1][11] ),
    .B(_01594_),
    .X(_03094_));
 sky130_fd_sc_hd__o21bai_2 _08174_ (.A1(_03093_),
    .A2(_03094_),
    .B1_N(_01110_),
    .Y(_03095_));
 sky130_fd_sc_hd__or2b_2 _08175_ (.A(\rvsingle.dp.rf.rf[3][11] ),
    .B_N(_01566_),
    .X(_03096_));
 sky130_fd_sc_hd__o211a_2 _08176_ (.A1(_01558_),
    .A2(\rvsingle.dp.rf.rf[2][11] ),
    .B1(_01880_),
    .C1(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__o21ai_2 _08177_ (.A1(_03095_),
    .A2(_03097_),
    .B1(_02364_),
    .Y(_03098_));
 sky130_fd_sc_hd__nor2_2 _08178_ (.A(_01545_),
    .B(\rvsingle.dp.rf.rf[12][11] ),
    .Y(_03099_));
 sky130_fd_sc_hd__o21ai_2 _08179_ (.A1(\rvsingle.dp.rf.rf[13][11] ),
    .A2(_02379_),
    .B1(_01542_),
    .Y(_03100_));
 sky130_fd_sc_hd__o21a_2 _08180_ (.A1(_01594_),
    .A2(\rvsingle.dp.rf.rf[14][11] ),
    .B1(_01489_),
    .X(_03101_));
 sky130_fd_sc_hd__o21ai_2 _08181_ (.A1(\rvsingle.dp.rf.rf[15][11] ),
    .A2(_01508_),
    .B1(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__o211ai_2 _08182_ (.A1(_03099_),
    .A2(_03100_),
    .B1(_02410_),
    .C1(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__nor2_2 _08183_ (.A(_01630_),
    .B(\rvsingle.dp.rf.rf[10][11] ),
    .Y(_03104_));
 sky130_fd_sc_hd__o21ai_2 _08184_ (.A1(\rvsingle.dp.rf.rf[11][11] ),
    .A2(_01860_),
    .B1(_01880_),
    .Y(_03105_));
 sky130_fd_sc_hd__or2_2 _08185_ (.A(_01096_),
    .B(\rvsingle.dp.rf.rf[8][11] ),
    .X(_03106_));
 sky130_fd_sc_hd__o211ai_2 _08186_ (.A1(\rvsingle.dp.rf.rf[9][11] ),
    .A2(_02379_),
    .B1(_01542_),
    .C1(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__o211ai_2 _08187_ (.A1(_03104_),
    .A2(_03105_),
    .B1(_02329_),
    .C1(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__nand3_2 _08188_ (.A(_03103_),
    .B(_03108_),
    .C(_01505_),
    .Y(_03109_));
 sky130_fd_sc_hd__o211ai_2 _08189_ (.A1(_03092_),
    .A2(_03098_),
    .B1(_01377_),
    .C1(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__o211ai_2 _08190_ (.A1(_01150_),
    .A2(_01139_),
    .B1(_03087_),
    .C1(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__o221ai_2 _08191_ (.A1(_02473_),
    .A2(_02318_),
    .B1(_01961_),
    .B2(_03111_),
    .C1(_01580_),
    .Y(_03112_));
 sky130_fd_sc_hd__mux4_2 _08192_ (.A0(\rvsingle.dp.rf.rf[4][11] ),
    .A1(\rvsingle.dp.rf.rf[5][11] ),
    .A2(\rvsingle.dp.rf.rf[6][11] ),
    .A3(\rvsingle.dp.rf.rf[7][11] ),
    .S0(_01426_),
    .S1(_01433_),
    .X(_03113_));
 sky130_fd_sc_hd__nor2_2 _08193_ (.A(_02093_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__mux4_2 _08194_ (.A0(\rvsingle.dp.rf.rf[0][11] ),
    .A1(\rvsingle.dp.rf.rf[1][11] ),
    .A2(\rvsingle.dp.rf.rf[2][11] ),
    .A3(\rvsingle.dp.rf.rf[3][11] ),
    .S0(_02450_),
    .S1(_01708_),
    .X(_03115_));
 sky130_fd_sc_hd__o21ai_2 _08195_ (.A1(_02302_),
    .A2(_03115_),
    .B1(_01699_),
    .Y(_03116_));
 sky130_fd_sc_hd__mux4_2 _08196_ (.A0(\rvsingle.dp.rf.rf[12][11] ),
    .A1(\rvsingle.dp.rf.rf[13][11] ),
    .A2(\rvsingle.dp.rf.rf[14][11] ),
    .A3(\rvsingle.dp.rf.rf[15][11] ),
    .S0(_01416_),
    .S1(_01300_),
    .X(_03117_));
 sky130_fd_sc_hd__nor2_2 _08197_ (.A(_01726_),
    .B(\rvsingle.dp.rf.rf[10][11] ),
    .Y(_03118_));
 sky130_fd_sc_hd__o21ai_2 _08198_ (.A1(\rvsingle.dp.rf.rf[11][11] ),
    .A2(_01295_),
    .B1(_01953_),
    .Y(_03119_));
 sky130_fd_sc_hd__or2_2 _08199_ (.A(_01828_),
    .B(\rvsingle.dp.rf.rf[8][11] ),
    .X(_03120_));
 sky130_fd_sc_hd__o211ai_2 _08200_ (.A1(\rvsingle.dp.rf.rf[9][11] ),
    .A2(_02303_),
    .B1(_01308_),
    .C1(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__o211ai_2 _08201_ (.A1(_03118_),
    .A2(_03119_),
    .B1(_02543_),
    .C1(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__o211ai_2 _08202_ (.A1(_01422_),
    .A2(_03117_),
    .B1(_03122_),
    .C1(_01221_),
    .Y(_03123_));
 sky130_fd_sc_hd__o211ai_2 _08203_ (.A1(_03114_),
    .A2(_03116_),
    .B1(_01315_),
    .C1(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__or2_2 _08204_ (.A(_01725_),
    .B(\rvsingle.dp.rf.rf[22][11] ),
    .X(_03125_));
 sky130_fd_sc_hd__o211a_2 _08205_ (.A1(_01295_),
    .A2(\rvsingle.dp.rf.rf[23][11] ),
    .B1(_01808_),
    .C1(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__or2_2 _08206_ (.A(_01191_),
    .B(\rvsingle.dp.rf.rf[20][11] ),
    .X(_03127_));
 sky130_fd_sc_hd__o211ai_2 _08207_ (.A1(\rvsingle.dp.rf.rf[21][11] ),
    .A2(_02303_),
    .B1(_01308_),
    .C1(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__nand2_2 _08208_ (.A(_03128_),
    .B(_02291_),
    .Y(_03129_));
 sky130_fd_sc_hd__mux4_2 _08209_ (.A0(\rvsingle.dp.rf.rf[16][11] ),
    .A1(\rvsingle.dp.rf.rf[17][11] ),
    .A2(\rvsingle.dp.rf.rf[18][11] ),
    .A3(\rvsingle.dp.rf.rf[19][11] ),
    .S0(_01416_),
    .S1(_01300_),
    .X(_03130_));
 sky130_fd_sc_hd__o22ai_2 _08210_ (.A1(_03126_),
    .A2(_03129_),
    .B1(_03130_),
    .B2(_01694_),
    .Y(_03131_));
 sky130_fd_sc_hd__mux4_2 _08211_ (.A0(\rvsingle.dp.rf.rf[28][11] ),
    .A1(\rvsingle.dp.rf.rf[29][11] ),
    .A2(\rvsingle.dp.rf.rf[30][11] ),
    .A3(\rvsingle.dp.rf.rf[31][11] ),
    .S0(_01730_),
    .S1(_01808_),
    .X(_03132_));
 sky130_fd_sc_hd__or2_2 _08212_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[24][11] ),
    .X(_03133_));
 sky130_fd_sc_hd__o211ai_2 _08213_ (.A1(\rvsingle.dp.rf.rf[25][11] ),
    .A2(_01827_),
    .B1(_01308_),
    .C1(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__or2_2 _08214_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[26][11] ),
    .X(_03135_));
 sky130_fd_sc_hd__o211ai_2 _08215_ (.A1(_02275_),
    .A2(\rvsingle.dp.rf.rf[27][11] ),
    .B1(_01433_),
    .C1(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__a31oi_2 _08216_ (.A1(_02543_),
    .A2(_03134_),
    .A3(_03136_),
    .B1(_01217_),
    .Y(_03137_));
 sky130_fd_sc_hd__o21ai_2 _08217_ (.A1(_02093_),
    .A2(_03132_),
    .B1(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__o211ai_2 _08218_ (.A1(_01447_),
    .A2(_03131_),
    .B1(_03138_),
    .C1(_02315_),
    .Y(_03139_));
 sky130_fd_sc_hd__o211a_2 _08219_ (.A1(_01201_),
    .A2(_01351_),
    .B1(_03124_),
    .C1(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__nand2_2 _08220_ (.A(_03112_),
    .B(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__o21a_2 _08221_ (.A1(_01483_),
    .A2(_02260_),
    .B1(_01177_),
    .X(_03142_));
 sky130_fd_sc_hd__a211oi_2 _08222_ (.A1(_03111_),
    .A2(_01870_),
    .B1(_01485_),
    .C1(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__mux4_2 _08223_ (.A0(\rvsingle.dp.rf.rf[20][10] ),
    .A1(\rvsingle.dp.rf.rf[21][10] ),
    .A2(\rvsingle.dp.rf.rf[22][10] ),
    .A3(\rvsingle.dp.rf.rf[23][10] ),
    .S0(_02176_),
    .S1(_01696_),
    .X(_03144_));
 sky130_fd_sc_hd__nor2_2 _08224_ (.A(_01422_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__mux4_2 _08225_ (.A0(\rvsingle.dp.rf.rf[16][10] ),
    .A1(\rvsingle.dp.rf.rf[17][10] ),
    .A2(\rvsingle.dp.rf.rf[18][10] ),
    .A3(\rvsingle.dp.rf.rf[19][10] ),
    .S0(_01328_),
    .S1(_01455_),
    .X(_03146_));
 sky130_fd_sc_hd__o21ai_2 _08226_ (.A1(_02302_),
    .A2(_03146_),
    .B1(_02447_),
    .Y(_03147_));
 sky130_fd_sc_hd__mux4_2 _08227_ (.A0(\rvsingle.dp.rf.rf[28][10] ),
    .A1(\rvsingle.dp.rf.rf[29][10] ),
    .A2(\rvsingle.dp.rf.rf[30][10] ),
    .A3(\rvsingle.dp.rf.rf[31][10] ),
    .S0(_02450_),
    .S1(_01708_),
    .X(_03148_));
 sky130_fd_sc_hd__mux2_2 _08228_ (.A0(\rvsingle.dp.rf.rf[24][10] ),
    .A1(\rvsingle.dp.rf.rf[25][10] ),
    .S(_01349_),
    .X(_03149_));
 sky130_fd_sc_hd__or2_2 _08229_ (.A(_01327_),
    .B(\rvsingle.dp.rf.rf[26][10] ),
    .X(_03150_));
 sky130_fd_sc_hd__o211a_2 _08230_ (.A1(_01294_),
    .A2(\rvsingle.dp.rf.rf[27][10] ),
    .B1(_01243_),
    .C1(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__a211o_2 _08231_ (.A1(_03149_),
    .A2(_02285_),
    .B1(_01444_),
    .C1(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__o211ai_2 _08232_ (.A1(_01422_),
    .A2(_03148_),
    .B1(_02438_),
    .C1(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__o211ai_2 _08233_ (.A1(_03145_),
    .A2(_03147_),
    .B1(_01187_),
    .C1(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__mux4_2 _08234_ (.A0(\rvsingle.dp.rf.rf[8][10] ),
    .A1(\rvsingle.dp.rf.rf[9][10] ),
    .A2(\rvsingle.dp.rf.rf[10][10] ),
    .A3(\rvsingle.dp.rf.rf[11][10] ),
    .S0(_02450_),
    .S1(_01708_),
    .X(_03155_));
 sky130_fd_sc_hd__or2_2 _08235_ (.A(_01725_),
    .B(\rvsingle.dp.rf.rf[12][10] ),
    .X(_03156_));
 sky130_fd_sc_hd__o211ai_2 _08236_ (.A1(\rvsingle.dp.rf.rf[13][10] ),
    .A2(_01901_),
    .B1(_02285_),
    .C1(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__o21a_2 _08237_ (.A1(_01903_),
    .A2(\rvsingle.dp.rf.rf[14][10] ),
    .B1(_01243_),
    .X(_03158_));
 sky130_fd_sc_hd__o21ai_2 _08238_ (.A1(\rvsingle.dp.rf.rf[15][10] ),
    .A2(_01901_),
    .B1(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__nand3_2 _08239_ (.A(_03157_),
    .B(_02291_),
    .C(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__o211ai_2 _08240_ (.A1(_02302_),
    .A2(_03155_),
    .B1(_03160_),
    .C1(_02438_),
    .Y(_03161_));
 sky130_fd_sc_hd__mux4_2 _08241_ (.A0(\rvsingle.dp.rf.rf[4][10] ),
    .A1(\rvsingle.dp.rf.rf[5][10] ),
    .A2(\rvsingle.dp.rf.rf[6][10] ),
    .A3(\rvsingle.dp.rf.rf[7][10] ),
    .S0(_01416_),
    .S1(_01708_),
    .X(_03162_));
 sky130_fd_sc_hd__nor2_2 _08242_ (.A(_01726_),
    .B(\rvsingle.dp.rf.rf[2][10] ),
    .Y(_03163_));
 sky130_fd_sc_hd__o21ai_2 _08243_ (.A1(\rvsingle.dp.rf.rf[3][10] ),
    .A2(_01827_),
    .B1(_01808_),
    .Y(_03164_));
 sky130_fd_sc_hd__or2_2 _08244_ (.A(_01191_),
    .B(\rvsingle.dp.rf.rf[0][10] ),
    .X(_03165_));
 sky130_fd_sc_hd__o211ai_2 _08245_ (.A1(\rvsingle.dp.rf.rf[1][10] ),
    .A2(_01295_),
    .B1(_01308_),
    .C1(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__o211ai_2 _08246_ (.A1(_03163_),
    .A2(_03164_),
    .B1(_02543_),
    .C1(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__o211ai_2 _08247_ (.A1(_01422_),
    .A2(_03162_),
    .B1(_03167_),
    .C1(_01699_),
    .Y(_03168_));
 sky130_fd_sc_hd__nand3_2 _08248_ (.A(_01315_),
    .B(_03161_),
    .C(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_2 _08249_ (.A(_03154_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__nand2_2 _08250_ (.A(_02375_),
    .B(Instr[30]),
    .Y(_03171_));
 sky130_fd_sc_hd__nor2_2 _08251_ (.A(_01619_),
    .B(\rvsingle.dp.rf.rf[10][10] ),
    .Y(_03172_));
 sky130_fd_sc_hd__o21ai_2 _08252_ (.A1(\rvsingle.dp.rf.rf[11][10] ),
    .A2(_01677_),
    .B1(_02320_),
    .Y(_03173_));
 sky130_fd_sc_hd__or2b_2 _08253_ (.A(\rvsingle.dp.rf.rf[9][10] ),
    .B_N(_01594_),
    .X(_03174_));
 sky130_fd_sc_hd__o211ai_2 _08254_ (.A1(_01595_),
    .A2(\rvsingle.dp.rf.rf[8][10] ),
    .B1(_03174_),
    .C1(_02485_),
    .Y(_03175_));
 sky130_fd_sc_hd__o211ai_2 _08255_ (.A1(_03172_),
    .A2(_03173_),
    .B1(_03175_),
    .C1(_01600_),
    .Y(_03176_));
 sky130_fd_sc_hd__nor2_2 _08256_ (.A(_01780_),
    .B(\rvsingle.dp.rf.rf[14][10] ),
    .Y(_03177_));
 sky130_fd_sc_hd__and2b_2 _08257_ (.A_N(\rvsingle.dp.rf.rf[15][10] ),
    .B(_01769_),
    .X(_03178_));
 sky130_fd_sc_hd__o21ba_2 _08258_ (.A1(_01136_),
    .A2(\rvsingle.dp.rf.rf[12][10] ),
    .B1_N(_01519_),
    .X(_03179_));
 sky130_fd_sc_hd__o21ai_2 _08259_ (.A1(_02478_),
    .A2(\rvsingle.dp.rf.rf[13][10] ),
    .B1(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__o311ai_2 _08260_ (.A1(_01092_),
    .A2(_03177_),
    .A3(_03178_),
    .B1(_01511_),
    .C1(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__nand3_2 _08261_ (.A(_03176_),
    .B(_02527_),
    .C(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__o21bai_2 _08262_ (.A1(_01763_),
    .A2(\rvsingle.dp.rf.rf[0][10] ),
    .B1_N(_01604_),
    .Y(_03183_));
 sky130_fd_sc_hd__and2b_2 _08263_ (.A_N(\rvsingle.dp.rf.rf[1][10] ),
    .B(_01743_),
    .X(_03184_));
 sky130_fd_sc_hd__o21ai_2 _08264_ (.A1(_03183_),
    .A2(_03184_),
    .B1(_02351_),
    .Y(_03185_));
 sky130_fd_sc_hd__or2b_2 _08265_ (.A(\rvsingle.dp.rf.rf[3][10] ),
    .B_N(_01561_),
    .X(_03186_));
 sky130_fd_sc_hd__o211a_2 _08266_ (.A1(_01518_),
    .A2(\rvsingle.dp.rf.rf[2][10] ),
    .B1(_02320_),
    .C1(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__nor2_2 _08267_ (.A(_01780_),
    .B(\rvsingle.dp.rf.rf[4][10] ),
    .Y(_03188_));
 sky130_fd_sc_hd__and2b_2 _08268_ (.A_N(\rvsingle.dp.rf.rf[5][10] ),
    .B(_02005_),
    .X(_03189_));
 sky130_fd_sc_hd__o21a_2 _08269_ (.A1(_01618_),
    .A2(\rvsingle.dp.rf.rf[6][10] ),
    .B1(_01551_),
    .X(_03190_));
 sky130_fd_sc_hd__o21ai_2 _08270_ (.A1(\rvsingle.dp.rf.rf[7][10] ),
    .A2(_02481_),
    .B1(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__o311ai_2 _08271_ (.A1(_01605_),
    .A2(_03188_),
    .A3(_03189_),
    .B1(_01511_),
    .C1(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__o211ai_2 _08272_ (.A1(_03185_),
    .A2(_03187_),
    .B1(_01156_),
    .C1(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand3_2 _08273_ (.A(_01593_),
    .B(_03182_),
    .C(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__nor2_2 _08274_ (.A(_01268_),
    .B(\rvsingle.dp.rf.rf[16][10] ),
    .Y(_03195_));
 sky130_fd_sc_hd__and2b_2 _08275_ (.A_N(\rvsingle.dp.rf.rf[17][10] ),
    .B(_01743_),
    .X(_03196_));
 sky130_fd_sc_hd__or2b_2 _08276_ (.A(\rvsingle.dp.rf.rf[19][10] ),
    .B_N(_01492_),
    .X(_03197_));
 sky130_fd_sc_hd__o211ai_2 _08277_ (.A1(_01268_),
    .A2(\rvsingle.dp.rf.rf[18][10] ),
    .B1(_02059_),
    .C1(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__o311ai_2 _08278_ (.A1(_01105_),
    .A2(_03195_),
    .A3(_03196_),
    .B1(_02483_),
    .C1(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__nor2_2 _08279_ (.A(_01268_),
    .B(\rvsingle.dp.rf.rf[22][10] ),
    .Y(_03200_));
 sky130_fd_sc_hd__and2b_2 _08280_ (.A_N(\rvsingle.dp.rf.rf[23][10] ),
    .B(_01743_),
    .X(_03201_));
 sky130_fd_sc_hd__o21ba_2 _08281_ (.A1(_01618_),
    .A2(\rvsingle.dp.rf.rf[20][10] ),
    .B1_N(_01489_),
    .X(_03202_));
 sky130_fd_sc_hd__o21ai_2 _08282_ (.A1(_02481_),
    .A2(\rvsingle.dp.rf.rf[21][10] ),
    .B1(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__o311ai_2 _08283_ (.A1(_01092_),
    .A2(_03200_),
    .A3(_03201_),
    .B1(_01511_),
    .C1(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__nand3_2 _08284_ (.A(_01853_),
    .B(_03199_),
    .C(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__o21bai_2 _08285_ (.A1(_01567_),
    .A2(\rvsingle.dp.rf.rf[24][10] ),
    .B1_N(_01604_),
    .Y(_03206_));
 sky130_fd_sc_hd__and2b_2 _08286_ (.A_N(\rvsingle.dp.rf.rf[25][10] ),
    .B(_01797_),
    .X(_03207_));
 sky130_fd_sc_hd__o21ai_2 _08287_ (.A1(_03206_),
    .A2(_03207_),
    .B1(_02483_),
    .Y(_03208_));
 sky130_fd_sc_hd__or2b_2 _08288_ (.A(\rvsingle.dp.rf.rf[27][10] ),
    .B_N(_01255_),
    .X(_03209_));
 sky130_fd_sc_hd__o211a_2 _08289_ (.A1(_01614_),
    .A2(\rvsingle.dp.rf.rf[26][10] ),
    .B1(_02320_),
    .C1(_03209_),
    .X(_03210_));
 sky130_fd_sc_hd__nor2_2 _08290_ (.A(_01878_),
    .B(\rvsingle.dp.rf.rf[28][10] ),
    .Y(_03211_));
 sky130_fd_sc_hd__and2b_2 _08291_ (.A_N(\rvsingle.dp.rf.rf[29][10] ),
    .B(_02005_),
    .X(_03212_));
 sky130_fd_sc_hd__or2b_2 _08292_ (.A(\rvsingle.dp.rf.rf[31][10] ),
    .B_N(_01267_),
    .X(_03213_));
 sky130_fd_sc_hd__o211ai_2 _08293_ (.A1(_01878_),
    .A2(\rvsingle.dp.rf.rf[30][10] ),
    .B1(_01520_),
    .C1(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__o311ai_2 _08294_ (.A1(_01605_),
    .A2(_03211_),
    .A3(_03212_),
    .B1(_01511_),
    .C1(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__o211ai_2 _08295_ (.A1(_03208_),
    .A2(_03210_),
    .B1(_02527_),
    .C1(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__nand3_2 _08296_ (.A(_03205_),
    .B(_01682_),
    .C(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__nand4_2 _08297_ (.A(_02505_),
    .B(_03194_),
    .C(_03217_),
    .D(_01083_),
    .Y(_03218_));
 sky130_fd_sc_hd__o211a_2 _08298_ (.A1(_02473_),
    .A2(_02318_),
    .B1(_03171_),
    .C1(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__a21oi_2 _08299_ (.A1(_03171_),
    .A2(_03218_),
    .B1(_01591_),
    .Y(_03220_));
 sky130_fd_sc_hd__o22ai_2 _08300_ (.A1(_02469_),
    .A2(_03170_),
    .B1(_03219_),
    .B2(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__and3_2 _08301_ (.A(_01246_),
    .B(_03154_),
    .C(_03169_),
    .X(_03222_));
 sky130_fd_sc_hd__o211ai_2 _08302_ (.A1(_01960_),
    .A2(_02102_),
    .B1(_03171_),
    .C1(_03218_),
    .Y(_03223_));
 sky130_fd_sc_hd__a31o_2 _08303_ (.A1(_01592_),
    .A2(_03194_),
    .A3(_03217_),
    .B1(_01178_),
    .X(_03224_));
 sky130_fd_sc_hd__or2_2 _08304_ (.A(Instr[30]),
    .B(_01481_),
    .X(_03225_));
 sky130_fd_sc_hd__nand3_2 _08305_ (.A(_03224_),
    .B(_03225_),
    .C(_01584_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand3_2 _08306_ (.A(_03222_),
    .B(_03223_),
    .C(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__nand2_2 _08307_ (.A(_03124_),
    .B(_03139_),
    .Y(_03228_));
 sky130_fd_sc_hd__o221a_2 _08308_ (.A1(_01065_),
    .A2(_01074_),
    .B1(_01961_),
    .B2(_03111_),
    .C1(_01580_),
    .X(_03229_));
 sky130_fd_sc_hd__o22ai_2 _08309_ (.A1(_02469_),
    .A2(_03228_),
    .B1(_03229_),
    .B2(_03143_),
    .Y(_03230_));
 sky130_fd_sc_hd__o2111ai_2 _08310_ (.A1(_03141_),
    .A2(_03143_),
    .B1(_03221_),
    .C1(_03227_),
    .D1(_03230_),
    .Y(_03231_));
 sky130_fd_sc_hd__inv_2 _08311_ (.A(Instr[28]),
    .Y(_03232_));
 sky130_fd_sc_hd__nor2_2 _08312_ (.A(_01513_),
    .B(\rvsingle.dp.rf.rf[14][8] ),
    .Y(_03233_));
 sky130_fd_sc_hd__o21ai_2 _08313_ (.A1(\rvsingle.dp.rf.rf[15][8] ),
    .A2(_01508_),
    .B1(_02059_),
    .Y(_03234_));
 sky130_fd_sc_hd__nor2_2 _08314_ (.A(_01493_),
    .B(\rvsingle.dp.rf.rf[12][8] ),
    .Y(_03235_));
 sky130_fd_sc_hd__o21ai_2 _08315_ (.A1(\rvsingle.dp.rf.rf[13][8] ),
    .A2(_01487_),
    .B1(_01496_),
    .Y(_03236_));
 sky130_fd_sc_hd__o221ai_2 _08316_ (.A1(_03233_),
    .A2(_03234_),
    .B1(_03235_),
    .B2(_03236_),
    .C1(_02488_),
    .Y(_03237_));
 sky130_fd_sc_hd__nor2_2 _08317_ (.A(_01878_),
    .B(\rvsingle.dp.rf.rf[8][8] ),
    .Y(_03238_));
 sky130_fd_sc_hd__o21ai_2 _08318_ (.A1(\rvsingle.dp.rf.rf[9][8] ),
    .A2(_01539_),
    .B1(_01542_),
    .Y(_03239_));
 sky130_fd_sc_hd__nor2_2 _08319_ (.A(_01499_),
    .B(\rvsingle.dp.rf.rf[10][8] ),
    .Y(_03240_));
 sky130_fd_sc_hd__o21ai_2 _08320_ (.A1(\rvsingle.dp.rf.rf[11][8] ),
    .A2(_01508_),
    .B1(_02059_),
    .Y(_03241_));
 sky130_fd_sc_hd__o221ai_2 _08321_ (.A1(_03238_),
    .A2(_03239_),
    .B1(_03240_),
    .B2(_03241_),
    .C1(_02483_),
    .Y(_03242_));
 sky130_fd_sc_hd__nand3_2 _08322_ (.A(_03237_),
    .B(_03242_),
    .C(_02527_),
    .Y(_03243_));
 sky130_fd_sc_hd__nor2_2 _08323_ (.A(_01137_),
    .B(\rvsingle.dp.rf.rf[2][8] ),
    .Y(_03244_));
 sky130_fd_sc_hd__o21ai_2 _08324_ (.A1(\rvsingle.dp.rf.rf[3][8] ),
    .A2(_02478_),
    .B1(_01523_),
    .Y(_03245_));
 sky130_fd_sc_hd__or2_2 _08325_ (.A(_02627_),
    .B(\rvsingle.dp.rf.rf[0][8] ),
    .X(_03246_));
 sky130_fd_sc_hd__o211ai_2 _08326_ (.A1(\rvsingle.dp.rf.rf[1][8] ),
    .A2(_02478_),
    .B1(_02395_),
    .C1(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__o211ai_2 _08327_ (.A1(_03244_),
    .A2(_03245_),
    .B1(_03247_),
    .C1(_02483_),
    .Y(_03248_));
 sky130_fd_sc_hd__nor2_2 _08328_ (.A(_01137_),
    .B(\rvsingle.dp.rf.rf[6][8] ),
    .Y(_03249_));
 sky130_fd_sc_hd__o21ai_2 _08329_ (.A1(\rvsingle.dp.rf.rf[7][8] ),
    .A2(_01487_),
    .B1(_01523_),
    .Y(_03250_));
 sky130_fd_sc_hd__or2_2 _08330_ (.A(_01267_),
    .B(\rvsingle.dp.rf.rf[4][8] ),
    .X(_03251_));
 sky130_fd_sc_hd__o211ai_2 _08331_ (.A1(\rvsingle.dp.rf.rf[5][8] ),
    .A2(_02481_),
    .B1(_01496_),
    .C1(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__o211ai_2 _08332_ (.A1(_03249_),
    .A2(_03250_),
    .B1(_02488_),
    .C1(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__nand3_2 _08333_ (.A(_01853_),
    .B(_03248_),
    .C(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand3_2 _08334_ (.A(_01593_),
    .B(_03243_),
    .C(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__nor2_2 _08335_ (.A(_01878_),
    .B(\rvsingle.dp.rf.rf[28][8] ),
    .Y(_03256_));
 sky130_fd_sc_hd__and2b_2 _08336_ (.A_N(\rvsingle.dp.rf.rf[29][8] ),
    .B(_01650_),
    .X(_03257_));
 sky130_fd_sc_hd__buf_1 _08337_ (.A(_01135_),
    .X(_03258_));
 sky130_fd_sc_hd__o21a_2 _08338_ (.A1(_03258_),
    .A2(\rvsingle.dp.rf.rf[30][8] ),
    .B1(_01604_),
    .X(_03259_));
 sky130_fd_sc_hd__o21ai_2 _08339_ (.A1(\rvsingle.dp.rf.rf[31][8] ),
    .A2(_01677_),
    .B1(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__o311a_2 _08340_ (.A1(_01605_),
    .A2(_03256_),
    .A3(_03257_),
    .B1(_01511_),
    .C1(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__inv_2 _08341_ (.A(\rvsingle.dp.rf.rf[25][8] ),
    .Y(_03262_));
 sky130_fd_sc_hd__o21bai_2 _08342_ (.A1(_01763_),
    .A2(\rvsingle.dp.rf.rf[24][8] ),
    .B1_N(_01604_),
    .Y(_03263_));
 sky130_fd_sc_hd__a21oi_2 _08343_ (.A1(_03262_),
    .A2(_01744_),
    .B1(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__o21ai_2 _08344_ (.A1(_01558_),
    .A2(\rvsingle.dp.rf.rf[26][8] ),
    .B1(_01777_),
    .Y(_03265_));
 sky130_fd_sc_hd__and2b_2 _08345_ (.A_N(\rvsingle.dp.rf.rf[27][8] ),
    .B(_01769_),
    .X(_03266_));
 sky130_fd_sc_hd__o21ai_2 _08346_ (.A1(_03265_),
    .A2(_03266_),
    .B1(_02351_),
    .Y(_03267_));
 sky130_fd_sc_hd__o21ai_2 _08347_ (.A1(_03264_),
    .A2(_03267_),
    .B1(_01505_),
    .Y(_03268_));
 sky130_fd_sc_hd__nor2_2 _08348_ (.A(_01763_),
    .B(\rvsingle.dp.rf.rf[16][8] ),
    .Y(_03269_));
 sky130_fd_sc_hd__and2b_2 _08349_ (.A_N(\rvsingle.dp.rf.rf[17][8] ),
    .B(_03258_),
    .X(_03270_));
 sky130_fd_sc_hd__or2b_2 _08350_ (.A(\rvsingle.dp.rf.rf[19][8] ),
    .B_N(_01877_),
    .X(_03271_));
 sky130_fd_sc_hd__o211ai_2 _08351_ (.A1(_01545_),
    .A2(\rvsingle.dp.rf.rf[18][8] ),
    .B1(_02031_),
    .C1(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__o311ai_2 _08352_ (.A1(_01531_),
    .A2(_03269_),
    .A3(_03270_),
    .B1(_01131_),
    .C1(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__nor2_2 _08353_ (.A(_01763_),
    .B(\rvsingle.dp.rf.rf[20][8] ),
    .Y(_03274_));
 sky130_fd_sc_hd__and2b_2 _08354_ (.A_N(\rvsingle.dp.rf.rf[21][8] ),
    .B(_03258_),
    .X(_03275_));
 sky130_fd_sc_hd__or2b_2 _08355_ (.A(\rvsingle.dp.rf.rf[23][8] ),
    .B_N(_01877_),
    .X(_03276_));
 sky130_fd_sc_hd__o211ai_2 _08356_ (.A1(_01545_),
    .A2(\rvsingle.dp.rf.rf[22][8] ),
    .B1(_02031_),
    .C1(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__o311ai_2 _08357_ (.A1(_01531_),
    .A2(_03274_),
    .A3(_03275_),
    .B1(_02410_),
    .C1(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__nand3_2 _08358_ (.A(_01853_),
    .B(_03273_),
    .C(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__o211ai_2 _08359_ (.A1(_03261_),
    .A2(_03268_),
    .B1(_01146_),
    .C1(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__nand4_2 _08360_ (.A(_03255_),
    .B(_01083_),
    .C(_02505_),
    .D(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__o21ai_2 _08361_ (.A1(_03232_),
    .A2(_01537_),
    .B1(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand2_2 _08362_ (.A(_03282_),
    .B(_01584_),
    .Y(_03283_));
 sky130_fd_sc_hd__mux2_2 _08363_ (.A0(\rvsingle.dp.rf.rf[4][8] ),
    .A1(\rvsingle.dp.rf.rf[5][8] ),
    .S(_01420_),
    .X(_03284_));
 sky130_fd_sc_hd__or2_2 _08364_ (.A(_01328_),
    .B(\rvsingle.dp.rf.rf[6][8] ),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_2 _08365_ (.A1(_01424_),
    .A2(\rvsingle.dp.rf.rf[7][8] ),
    .B1(_01244_),
    .C1(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__a211oi_2 _08366_ (.A1(_03284_),
    .A2(_01309_),
    .B1(_01422_),
    .C1(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__mux4_2 _08367_ (.A0(\rvsingle.dp.rf.rf[0][8] ),
    .A1(\rvsingle.dp.rf.rf[1][8] ),
    .A2(\rvsingle.dp.rf.rf[2][8] ),
    .A3(\rvsingle.dp.rf.rf[3][8] ),
    .S0(_01730_),
    .S1(_01808_),
    .X(_03288_));
 sky130_fd_sc_hd__o21ai_2 _08368_ (.A1(_01694_),
    .A2(_03288_),
    .B1(_01699_),
    .Y(_03289_));
 sky130_fd_sc_hd__mux4_2 _08369_ (.A0(\rvsingle.dp.rf.rf[12][8] ),
    .A1(\rvsingle.dp.rf.rf[13][8] ),
    .A2(\rvsingle.dp.rf.rf[14][8] ),
    .A3(\rvsingle.dp.rf.rf[15][8] ),
    .S0(_01241_),
    .S1(_01953_),
    .X(_03290_));
 sky130_fd_sc_hd__nor2_2 _08370_ (.A(_01329_),
    .B(\rvsingle.dp.rf.rf[8][8] ),
    .Y(_03291_));
 sky130_fd_sc_hd__o21ai_2 _08371_ (.A1(\rvsingle.dp.rf.rf[9][8] ),
    .A2(_01424_),
    .B1(_01716_),
    .Y(_03292_));
 sky130_fd_sc_hd__o21a_2 _08372_ (.A1(_01426_),
    .A2(\rvsingle.dp.rf.rf[10][8] ),
    .B1(_01427_),
    .X(_03293_));
 sky130_fd_sc_hd__o21ai_2 _08373_ (.A1(\rvsingle.dp.rf.rf[11][8] ),
    .A2(_01424_),
    .B1(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__o211ai_2 _08374_ (.A1(_03291_),
    .A2(_03292_),
    .B1(_01721_),
    .C1(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__o211ai_2 _08375_ (.A1(_02093_),
    .A2(_03290_),
    .B1(_03295_),
    .C1(_01447_),
    .Y(_03296_));
 sky130_fd_sc_hd__o21ai_2 _08376_ (.A1(_03287_),
    .A2(_03289_),
    .B1(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__mux2_2 _08377_ (.A0(\rvsingle.dp.rf.rf[26][8] ),
    .A1(\rvsingle.dp.rf.rf[27][8] ),
    .S(_01707_),
    .X(_03298_));
 sky130_fd_sc_hd__or2_2 _08378_ (.A(_02440_),
    .B(\rvsingle.dp.rf.rf[24][8] ),
    .X(_03299_));
 sky130_fd_sc_hd__o211a_2 _08379_ (.A1(\rvsingle.dp.rf.rf[25][8] ),
    .A2(_01901_),
    .B1(_02285_),
    .C1(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__a211oi_2 _08380_ (.A1(_01200_),
    .A2(_03298_),
    .B1(_03300_),
    .C1(_01694_),
    .Y(_03301_));
 sky130_fd_sc_hd__mux4_2 _08381_ (.A0(\rvsingle.dp.rf.rf[28][8] ),
    .A1(\rvsingle.dp.rf.rf[29][8] ),
    .A2(\rvsingle.dp.rf.rf[30][8] ),
    .A3(\rvsingle.dp.rf.rf[31][8] ),
    .S0(_01730_),
    .S1(_01953_),
    .X(_03302_));
 sky130_fd_sc_hd__o21ai_2 _08382_ (.A1(_02093_),
    .A2(_03302_),
    .B1(_01221_),
    .Y(_03303_));
 sky130_fd_sc_hd__mux4_2 _08383_ (.A0(\rvsingle.dp.rf.rf[16][8] ),
    .A1(\rvsingle.dp.rf.rf[17][8] ),
    .A2(\rvsingle.dp.rf.rf[18][8] ),
    .A3(\rvsingle.dp.rf.rf[19][8] ),
    .S0(_01730_),
    .S1(_01808_),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_2 _08384_ (.A0(\rvsingle.dp.rf.rf[20][8] ),
    .A1(\rvsingle.dp.rf.rf[21][8] ),
    .S(_01191_),
    .X(_03305_));
 sky130_fd_sc_hd__o21a_2 _08385_ (.A1(_01240_),
    .A2(\rvsingle.dp.rf.rf[22][8] ),
    .B1(_01454_),
    .X(_03306_));
 sky130_fd_sc_hd__o21a_2 _08386_ (.A1(_02929_),
    .A2(\rvsingle.dp.rf.rf[23][8] ),
    .B1(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__a211o_2 _08387_ (.A1(_03305_),
    .A2(_01716_),
    .B1(_01460_),
    .C1(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__o211ai_2 _08388_ (.A1(_01694_),
    .A2(_03304_),
    .B1(_03308_),
    .C1(_01699_),
    .Y(_03309_));
 sky130_fd_sc_hd__o211ai_2 _08389_ (.A1(_03301_),
    .A2(_03303_),
    .B1(_03309_),
    .C1(_02315_),
    .Y(_03310_));
 sky130_fd_sc_hd__o211a_2 _08390_ (.A1(_01188_),
    .A2(_03297_),
    .B1(_03310_),
    .C1(_01247_),
    .X(_03311_));
 sky130_fd_sc_hd__o221ai_2 _08391_ (.A1(_01960_),
    .A2(_02102_),
    .B1(_01084_),
    .B2(_03232_),
    .C1(_03281_),
    .Y(_03312_));
 sky130_fd_sc_hd__nand3_2 _08392_ (.A(_03283_),
    .B(_03311_),
    .C(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__o221a_2 _08393_ (.A1(_01960_),
    .A2(_02102_),
    .B1(_01084_),
    .B2(_03232_),
    .C1(_03281_),
    .X(_03314_));
 sky130_fd_sc_hd__nand2_2 _08394_ (.A(_01961_),
    .B(Instr[28]),
    .Y(_03315_));
 sky130_fd_sc_hd__a21oi_2 _08395_ (.A1(_03315_),
    .A2(_03281_),
    .B1(_01486_),
    .Y(_03316_));
 sky130_fd_sc_hd__o21bai_2 _08396_ (.A1(_03314_),
    .A2(_03316_),
    .B1_N(_03311_),
    .Y(_03317_));
 sky130_fd_sc_hd__nand2_2 _08397_ (.A(_01178_),
    .B(Instr[29]),
    .Y(_03318_));
 sky130_fd_sc_hd__o21bai_2 _08398_ (.A1(_02030_),
    .A2(\rvsingle.dp.rf.rf[8][9] ),
    .B1_N(_01104_),
    .Y(_03319_));
 sky130_fd_sc_hd__and2b_2 _08399_ (.A_N(\rvsingle.dp.rf.rf[9][9] ),
    .B(_01607_),
    .X(_03320_));
 sky130_fd_sc_hd__o21ai_2 _08400_ (.A1(_03319_),
    .A2(_03320_),
    .B1(_02483_),
    .Y(_03321_));
 sky130_fd_sc_hd__or2b_2 _08401_ (.A(\rvsingle.dp.rf.rf[11][9] ),
    .B_N(_03258_),
    .X(_03322_));
 sky130_fd_sc_hd__o211a_2 _08402_ (.A1(_01562_),
    .A2(\rvsingle.dp.rf.rf[10][9] ),
    .B1(_01620_),
    .C1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__nor2_2 _08403_ (.A(_01268_),
    .B(\rvsingle.dp.rf.rf[12][9] ),
    .Y(_03324_));
 sky130_fd_sc_hd__and2b_2 _08404_ (.A_N(\rvsingle.dp.rf.rf[13][9] ),
    .B(_01743_),
    .X(_03325_));
 sky130_fd_sc_hd__or2b_2 _08405_ (.A(\rvsingle.dp.rf.rf[15][9] ),
    .B_N(_01492_),
    .X(_03326_));
 sky130_fd_sc_hd__o211ai_2 _08406_ (.A1(_01268_),
    .A2(\rvsingle.dp.rf.rf[14][9] ),
    .B1(_02059_),
    .C1(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__o311ai_2 _08407_ (.A1(_01105_),
    .A2(_03324_),
    .A3(_03325_),
    .B1(_01511_),
    .C1(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__o211ai_2 _08408_ (.A1(_03321_),
    .A2(_03323_),
    .B1(_02527_),
    .C1(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__nor2_2 _08409_ (.A(_01268_),
    .B(\rvsingle.dp.rf.rf[0][9] ),
    .Y(_03330_));
 sky130_fd_sc_hd__and2b_2 _08410_ (.A_N(\rvsingle.dp.rf.rf[1][9] ),
    .B(_01743_),
    .X(_03331_));
 sky130_fd_sc_hd__or2b_2 _08411_ (.A(\rvsingle.dp.rf.rf[3][9] ),
    .B_N(_01492_),
    .X(_03332_));
 sky130_fd_sc_hd__o211ai_2 _08412_ (.A1(_01513_),
    .A2(\rvsingle.dp.rf.rf[2][9] ),
    .B1(_02059_),
    .C1(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__o311ai_2 _08413_ (.A1(_01105_),
    .A2(_03330_),
    .A3(_03331_),
    .B1(_02483_),
    .C1(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__nor2_2 _08414_ (.A(_01268_),
    .B(\rvsingle.dp.rf.rf[4][9] ),
    .Y(_03335_));
 sky130_fd_sc_hd__and2b_2 _08415_ (.A_N(\rvsingle.dp.rf.rf[5][9] ),
    .B(_01743_),
    .X(_03336_));
 sky130_fd_sc_hd__or2b_2 _08416_ (.A(\rvsingle.dp.rf.rf[7][9] ),
    .B_N(_01492_),
    .X(_03337_));
 sky130_fd_sc_hd__o211ai_2 _08417_ (.A1(_01513_),
    .A2(\rvsingle.dp.rf.rf[6][9] ),
    .B1(_01490_),
    .C1(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__o311ai_2 _08418_ (.A1(_01105_),
    .A2(_03335_),
    .A3(_03336_),
    .B1(_02488_),
    .C1(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__nand3_2 _08419_ (.A(_01634_),
    .B(_03334_),
    .C(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__nand3_2 _08420_ (.A(_01593_),
    .B(_03329_),
    .C(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__nor2_2 _08421_ (.A(_01603_),
    .B(\rvsingle.dp.rf.rf[30][9] ),
    .Y(_03342_));
 sky130_fd_sc_hd__o21ai_2 _08422_ (.A1(\rvsingle.dp.rf.rf[31][9] ),
    .A2(_01796_),
    .B1(_01660_),
    .Y(_03343_));
 sky130_fd_sc_hd__or2b_2 _08423_ (.A(\rvsingle.dp.rf.rf[29][9] ),
    .B_N(_01618_),
    .X(_03344_));
 sky130_fd_sc_hd__o211ai_2 _08424_ (.A1(_01562_),
    .A2(\rvsingle.dp.rf.rf[28][9] ),
    .B1(_03344_),
    .C1(_02485_),
    .Y(_03345_));
 sky130_fd_sc_hd__o211ai_2 _08425_ (.A1(_03342_),
    .A2(_03343_),
    .B1(_03345_),
    .C1(_01632_),
    .Y(_03346_));
 sky130_fd_sc_hd__o21a_2 _08426_ (.A1(_02005_),
    .A2(\rvsingle.dp.rf.rf[26][9] ),
    .B1(_01104_),
    .X(_03347_));
 sky130_fd_sc_hd__o21ai_2 _08427_ (.A1(\rvsingle.dp.rf.rf[27][9] ),
    .A2(_01796_),
    .B1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__o21ba_2 _08428_ (.A1(_02005_),
    .A2(\rvsingle.dp.rf.rf[24][9] ),
    .B1_N(_01530_),
    .X(_03349_));
 sky130_fd_sc_hd__o21ai_2 _08429_ (.A1(_01796_),
    .A2(\rvsingle.dp.rf.rf[25][9] ),
    .B1(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__nand3_2 _08430_ (.A(_01768_),
    .B(_03348_),
    .C(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__nand3_2 _08431_ (.A(_03346_),
    .B(_03351_),
    .C(_01116_),
    .Y(_03352_));
 sky130_fd_sc_hd__o21bai_2 _08432_ (.A1(_02030_),
    .A2(\rvsingle.dp.rf.rf[16][9] ),
    .B1_N(_01104_),
    .Y(_03353_));
 sky130_fd_sc_hd__and2b_2 _08433_ (.A_N(\rvsingle.dp.rf.rf[17][9] ),
    .B(_01607_),
    .X(_03354_));
 sky130_fd_sc_hd__o21ai_2 _08434_ (.A1(_03353_),
    .A2(_03354_),
    .B1(_02483_),
    .Y(_03355_));
 sky130_fd_sc_hd__or2b_2 _08435_ (.A(\rvsingle.dp.rf.rf[19][9] ),
    .B_N(_03258_),
    .X(_03356_));
 sky130_fd_sc_hd__o211a_2 _08436_ (.A1(_01619_),
    .A2(\rvsingle.dp.rf.rf[18][9] ),
    .B1(_01620_),
    .C1(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__nor2_2 _08437_ (.A(_01499_),
    .B(\rvsingle.dp.rf.rf[20][9] ),
    .Y(_03358_));
 sky130_fd_sc_hd__and2b_2 _08438_ (.A_N(\rvsingle.dp.rf.rf[21][9] ),
    .B(_01125_),
    .X(_03359_));
 sky130_fd_sc_hd__or2b_2 _08439_ (.A(\rvsingle.dp.rf.rf[23][9] ),
    .B_N(_01492_),
    .X(_03360_));
 sky130_fd_sc_hd__o211ai_2 _08440_ (.A1(_01268_),
    .A2(\rvsingle.dp.rf.rf[22][9] ),
    .B1(_02059_),
    .C1(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__o311ai_2 _08441_ (.A1(_01605_),
    .A2(_03358_),
    .A3(_03359_),
    .B1(_01511_),
    .C1(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__o211ai_2 _08442_ (.A1(_03355_),
    .A2(_03357_),
    .B1(_01853_),
    .C1(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__nand3_2 _08443_ (.A(_03352_),
    .B(_03363_),
    .C(_01682_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand4_2 _08444_ (.A(_03341_),
    .B(_01481_),
    .C(_01592_),
    .D(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__o211a_2 _08445_ (.A1(_01960_),
    .A2(_02102_),
    .B1(_03318_),
    .C1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__a21oi_2 _08446_ (.A1(_03318_),
    .A2(_03365_),
    .B1(_01486_),
    .Y(_03367_));
 sky130_fd_sc_hd__mux4_2 _08447_ (.A0(\rvsingle.dp.rf.rf[8][9] ),
    .A1(\rvsingle.dp.rf.rf[9][9] ),
    .A2(\rvsingle.dp.rf.rf[10][9] ),
    .A3(\rvsingle.dp.rf.rf[11][9] ),
    .S0(_02176_),
    .S1(_01696_),
    .X(_03368_));
 sky130_fd_sc_hd__or2_2 _08448_ (.A(_01349_),
    .B(\rvsingle.dp.rf.rf[12][9] ),
    .X(_03369_));
 sky130_fd_sc_hd__o211ai_2 _08449_ (.A1(\rvsingle.dp.rf.rf[13][9] ),
    .A2(_02288_),
    .B1(_01436_),
    .C1(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__o21a_2 _08450_ (.A1(_01468_),
    .A2(\rvsingle.dp.rf.rf[14][9] ),
    .B1(_01198_),
    .X(_03371_));
 sky130_fd_sc_hd__o21ai_2 _08451_ (.A1(\rvsingle.dp.rf.rf[15][9] ),
    .A2(_01827_),
    .B1(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__a31oi_2 _08452_ (.A1(_03370_),
    .A2(_02291_),
    .A3(_03372_),
    .B1(_01217_),
    .Y(_03373_));
 sky130_fd_sc_hd__o21ai_2 _08453_ (.A1(_01711_),
    .A2(_03368_),
    .B1(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__mux4_2 _08454_ (.A0(\rvsingle.dp.rf.rf[0][9] ),
    .A1(\rvsingle.dp.rf.rf[1][9] ),
    .A2(\rvsingle.dp.rf.rf[2][9] ),
    .A3(\rvsingle.dp.rf.rf[3][9] ),
    .S0(_02176_),
    .S1(_02162_),
    .X(_03375_));
 sky130_fd_sc_hd__or2_2 _08455_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[4][9] ),
    .X(_03376_));
 sky130_fd_sc_hd__o211ai_2 _08456_ (.A1(\rvsingle.dp.rf.rf[5][9] ),
    .A2(_01827_),
    .B1(_01308_),
    .C1(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__o21a_2 _08457_ (.A1(_01468_),
    .A2(\rvsingle.dp.rf.rf[6][9] ),
    .B1(_01198_),
    .X(_03378_));
 sky130_fd_sc_hd__o21ai_2 _08458_ (.A1(\rvsingle.dp.rf.rf[7][9] ),
    .A2(_01295_),
    .B1(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__a31oi_2 _08459_ (.A1(_03377_),
    .A2(_02291_),
    .A3(_03379_),
    .B1(_01446_),
    .Y(_03380_));
 sky130_fd_sc_hd__o21ai_2 _08460_ (.A1(_01711_),
    .A2(_03375_),
    .B1(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__nand3_2 _08461_ (.A(_01315_),
    .B(_03374_),
    .C(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__mux4_2 _08462_ (.A0(\rvsingle.dp.rf.rf[28][9] ),
    .A1(\rvsingle.dp.rf.rf[29][9] ),
    .A2(\rvsingle.dp.rf.rf[30][9] ),
    .A3(\rvsingle.dp.rf.rf[31][9] ),
    .S0(_01426_),
    .S1(_01433_),
    .X(_03383_));
 sky130_fd_sc_hd__o21a_2 _08463_ (.A1(_02440_),
    .A2(\rvsingle.dp.rf.rf[26][9] ),
    .B1(_01243_),
    .X(_03384_));
 sky130_fd_sc_hd__o21ai_2 _08464_ (.A1(\rvsingle.dp.rf.rf[27][9] ),
    .A2(_02303_),
    .B1(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__or2_2 _08465_ (.A(_01349_),
    .B(\rvsingle.dp.rf.rf[24][9] ),
    .X(_03386_));
 sky130_fd_sc_hd__o211ai_2 _08466_ (.A1(\rvsingle.dp.rf.rf[25][9] ),
    .A2(_02288_),
    .B1(_01436_),
    .C1(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__a31oi_2 _08467_ (.A1(_02543_),
    .A2(_03385_),
    .A3(_03387_),
    .B1(_01217_),
    .Y(_03388_));
 sky130_fd_sc_hd__o21ai_2 _08468_ (.A1(_02093_),
    .A2(_03383_),
    .B1(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__mux4_2 _08469_ (.A0(\rvsingle.dp.rf.rf[20][9] ),
    .A1(\rvsingle.dp.rf.rf[21][9] ),
    .A2(\rvsingle.dp.rf.rf[22][9] ),
    .A3(\rvsingle.dp.rf.rf[23][9] ),
    .S0(_01328_),
    .S1(_01455_),
    .X(_03390_));
 sky130_fd_sc_hd__nor2_2 _08470_ (.A(\rvsingle.dp.rf.rf[19][9] ),
    .B(_02303_),
    .Y(_03391_));
 sky130_fd_sc_hd__o21ai_2 _08471_ (.A1(_01695_),
    .A2(\rvsingle.dp.rf.rf[18][9] ),
    .B1(_01433_),
    .Y(_03392_));
 sky130_fd_sc_hd__or2_2 _08472_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[16][9] ),
    .X(_03393_));
 sky130_fd_sc_hd__o211ai_2 _08473_ (.A1(\rvsingle.dp.rf.rf[17][9] ),
    .A2(_01827_),
    .B1(_01308_),
    .C1(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__o211ai_2 _08474_ (.A1(_03391_),
    .A2(_03392_),
    .B1(_02543_),
    .C1(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__o211ai_2 _08475_ (.A1(_01207_),
    .A2(_03390_),
    .B1(_03395_),
    .C1(_02447_),
    .Y(_03396_));
 sky130_fd_sc_hd__nand3_2 _08476_ (.A(_03389_),
    .B(_03396_),
    .C(_02315_),
    .Y(_03397_));
 sky130_fd_sc_hd__o211ai_2 _08477_ (.A1(_01351_),
    .A2(_01202_),
    .B1(_03382_),
    .C1(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__o21ai_2 _08478_ (.A1(_03366_),
    .A2(_03367_),
    .B1(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__a31o_2 _08479_ (.A1(_02505_),
    .A2(_03341_),
    .A3(_03364_),
    .B1(_02375_),
    .X(_03400_));
 sky130_fd_sc_hd__or2_2 _08480_ (.A(Instr[29]),
    .B(_01083_),
    .X(_03401_));
 sky130_fd_sc_hd__nand3_2 _08481_ (.A(_03400_),
    .B(_03401_),
    .C(_01584_),
    .Y(_03402_));
 sky130_fd_sc_hd__and3_2 _08482_ (.A(_01247_),
    .B(_03397_),
    .C(_03382_),
    .X(_03403_));
 sky130_fd_sc_hd__o211ai_2 _08483_ (.A1(_01960_),
    .A2(_02102_),
    .B1(_03318_),
    .C1(_03365_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand3_2 _08484_ (.A(_03402_),
    .B(_03403_),
    .C(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand4_2 _08485_ (.A(_03313_),
    .B(_03317_),
    .C(_03399_),
    .D(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__or2b_2 _08486_ (.A(\rvsingle.dp.rf.rf[27][13] ),
    .B_N(_01381_),
    .X(_03407_));
 sky130_fd_sc_hd__o211a_2 _08487_ (.A1(_01658_),
    .A2(\rvsingle.dp.rf.rf[26][13] ),
    .B1(_01880_),
    .C1(_03407_),
    .X(_03408_));
 sky130_fd_sc_hd__o21bai_2 _08488_ (.A1(_01607_),
    .A2(\rvsingle.dp.rf.rf[24][13] ),
    .B1_N(_01489_),
    .Y(_03409_));
 sky130_fd_sc_hd__and2b_2 _08489_ (.A_N(\rvsingle.dp.rf.rf[25][13] ),
    .B(_01136_),
    .X(_03410_));
 sky130_fd_sc_hd__o21ai_2 _08490_ (.A1(_03409_),
    .A2(_03410_),
    .B1(_02329_),
    .Y(_03411_));
 sky130_fd_sc_hd__nor2_2 _08491_ (.A(_01862_),
    .B(\rvsingle.dp.rf.rf[30][13] ),
    .Y(_03412_));
 sky130_fd_sc_hd__o21ai_2 _08492_ (.A1(\rvsingle.dp.rf.rf[31][13] ),
    .A2(_01087_),
    .B1(_01880_),
    .Y(_03413_));
 sky130_fd_sc_hd__o21ba_2 _08493_ (.A1(_01544_),
    .A2(\rvsingle.dp.rf.rf[28][13] ),
    .B1_N(_01610_),
    .X(_03414_));
 sky130_fd_sc_hd__o21ai_2 _08494_ (.A1(_01860_),
    .A2(\rvsingle.dp.rf.rf[29][13] ),
    .B1(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__o211ai_2 _08495_ (.A1(_03412_),
    .A2(_03413_),
    .B1(_03415_),
    .C1(_02323_),
    .Y(_03416_));
 sky130_fd_sc_hd__o211ai_2 _08496_ (.A1(_03408_),
    .A2(_03411_),
    .B1(_02491_),
    .C1(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__o21bai_2 _08497_ (.A1(_01769_),
    .A2(\rvsingle.dp.rf.rf[16][13] ),
    .B1_N(_01519_),
    .Y(_03418_));
 sky130_fd_sc_hd__and2b_2 _08498_ (.A_N(\rvsingle.dp.rf.rf[17][13] ),
    .B(_01498_),
    .X(_03419_));
 sky130_fd_sc_hd__o21ai_2 _08499_ (.A1(_03418_),
    .A2(_03419_),
    .B1(_01564_),
    .Y(_03420_));
 sky130_fd_sc_hd__or2b_2 _08500_ (.A(\rvsingle.dp.rf.rf[19][13] ),
    .B_N(_01381_),
    .X(_03421_));
 sky130_fd_sc_hd__o211a_2 _08501_ (.A1(_01097_),
    .A2(\rvsingle.dp.rf.rf[18][13] ),
    .B1(_01654_),
    .C1(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__o21ba_2 _08502_ (.A1(_01779_),
    .A2(\rvsingle.dp.rf.rf[20][13] ),
    .B1_N(_01610_),
    .X(_03423_));
 sky130_fd_sc_hd__o21ai_2 _08503_ (.A1(_02379_),
    .A2(\rvsingle.dp.rf.rf[21][13] ),
    .B1(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__o21a_2 _08504_ (.A1(_01544_),
    .A2(\rvsingle.dp.rf.rf[22][13] ),
    .B1(_01258_),
    .X(_03425_));
 sky130_fd_sc_hd__o21ai_2 _08505_ (.A1(\rvsingle.dp.rf.rf[23][13] ),
    .A2(_01860_),
    .B1(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand3_2 _08506_ (.A(_03424_),
    .B(_01111_),
    .C(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__o211ai_2 _08507_ (.A1(_03420_),
    .A2(_03422_),
    .B1(_02364_),
    .C1(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__nand3_2 _08508_ (.A(_03417_),
    .B(_03428_),
    .C(_01145_),
    .Y(_03429_));
 sky130_fd_sc_hd__nor2_2 _08509_ (.A(_01382_),
    .B(\rvsingle.dp.rf.rf[10][13] ),
    .Y(_03430_));
 sky130_fd_sc_hd__o21ai_2 _08510_ (.A1(\rvsingle.dp.rf.rf[11][13] ),
    .A2(_01860_),
    .B1(_01259_),
    .Y(_03431_));
 sky130_fd_sc_hd__or2b_2 _08511_ (.A(\rvsingle.dp.rf.rf[9][13] ),
    .B_N(_01096_),
    .X(_03432_));
 sky130_fd_sc_hd__o211ai_2 _08512_ (.A1(_02117_),
    .A2(\rvsingle.dp.rf.rf[8][13] ),
    .B1(_03432_),
    .C1(_01542_),
    .Y(_03433_));
 sky130_fd_sc_hd__o211ai_2 _08513_ (.A1(_03430_),
    .A2(_03431_),
    .B1(_03433_),
    .C1(_01131_),
    .Y(_03434_));
 sky130_fd_sc_hd__nor2_2 _08514_ (.A(_01607_),
    .B(\rvsingle.dp.rf.rf[14][13] ),
    .Y(_03435_));
 sky130_fd_sc_hd__and2b_2 _08515_ (.A_N(\rvsingle.dp.rf.rf[15][13] ),
    .B(_02627_),
    .X(_03436_));
 sky130_fd_sc_hd__o21ba_2 _08516_ (.A1(_01557_),
    .A2(\rvsingle.dp.rf.rf[12][13] ),
    .B1_N(_01103_),
    .X(_03437_));
 sky130_fd_sc_hd__o21ai_2 _08517_ (.A1(_01087_),
    .A2(\rvsingle.dp.rf.rf[13][13] ),
    .B1(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__o311ai_2 _08518_ (.A1(_02395_),
    .A2(_03435_),
    .A3(_03436_),
    .B1(_01502_),
    .C1(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand3_2 _08519_ (.A(_03434_),
    .B(_02491_),
    .C(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__nor2_2 _08520_ (.A(_01642_),
    .B(\rvsingle.dp.rf.rf[0][13] ),
    .Y(_03441_));
 sky130_fd_sc_hd__and2b_2 _08521_ (.A_N(\rvsingle.dp.rf.rf[1][13] ),
    .B(_01498_),
    .X(_03442_));
 sky130_fd_sc_hd__or2b_2 _08522_ (.A(\rvsingle.dp.rf.rf[3][13] ),
    .B_N(_01752_),
    .X(_03443_));
 sky130_fd_sc_hd__o211ai_2 _08523_ (.A1(_01642_),
    .A2(\rvsingle.dp.rf.rf[2][13] ),
    .B1(_01596_),
    .C1(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__o311ai_2 _08524_ (.A1(_01520_),
    .A2(_03441_),
    .A3(_03442_),
    .B1(_01564_),
    .C1(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__nor2_2 _08525_ (.A(_01642_),
    .B(\rvsingle.dp.rf.rf[4][13] ),
    .Y(_03446_));
 sky130_fd_sc_hd__and2b_2 _08526_ (.A_N(\rvsingle.dp.rf.rf[5][13] ),
    .B(_01498_),
    .X(_03447_));
 sky130_fd_sc_hd__or2b_2 _08527_ (.A(\rvsingle.dp.rf.rf[7][13] ),
    .B_N(_01752_),
    .X(_03448_));
 sky130_fd_sc_hd__o211ai_2 _08528_ (.A1(_01753_),
    .A2(\rvsingle.dp.rf.rf[6][13] ),
    .B1(_01596_),
    .C1(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__o311ai_2 _08529_ (.A1(_01520_),
    .A2(_03446_),
    .A3(_03447_),
    .B1(_01502_),
    .C1(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__nand3_2 _08530_ (.A(_01156_),
    .B(_03445_),
    .C(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand3_2 _08531_ (.A(_01377_),
    .B(_03440_),
    .C(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__o211ai_2 _08532_ (.A1(_01150_),
    .A2(_01139_),
    .B1(_03429_),
    .C1(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__a211oi_2 _08533_ (.A1(_03453_),
    .A2(_01870_),
    .B1(_01485_),
    .C1(_03142_),
    .Y(_03454_));
 sky130_fd_sc_hd__a21oi_2 _08534_ (.A1(_03453_),
    .A2(_01084_),
    .B1(_03142_),
    .Y(_03455_));
 sky130_fd_sc_hd__mux4_2 _08535_ (.A0(\rvsingle.dp.rf.rf[16][13] ),
    .A1(\rvsingle.dp.rf.rf[17][13] ),
    .A2(\rvsingle.dp.rf.rf[18][13] ),
    .A3(\rvsingle.dp.rf.rf[19][13] ),
    .S0(_01416_),
    .S1(_01696_),
    .X(_03456_));
 sky130_fd_sc_hd__nor2_2 _08536_ (.A(_01711_),
    .B(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__mux4_2 _08537_ (.A0(\rvsingle.dp.rf.rf[20][13] ),
    .A1(\rvsingle.dp.rf.rf[21][13] ),
    .A2(\rvsingle.dp.rf.rf[22][13] ),
    .A3(\rvsingle.dp.rf.rf[23][13] ),
    .S0(_01328_),
    .S1(_01470_),
    .X(_03458_));
 sky130_fd_sc_hd__o21ai_2 _08538_ (.A1(_01207_),
    .A2(_03458_),
    .B1(_02447_),
    .Y(_03459_));
 sky130_fd_sc_hd__mux4_2 _08539_ (.A0(\rvsingle.dp.rf.rf[24][13] ),
    .A1(\rvsingle.dp.rf.rf[25][13] ),
    .A2(\rvsingle.dp.rf.rf[26][13] ),
    .A3(\rvsingle.dp.rf.rf[27][13] ),
    .S0(_01468_),
    .S1(_01727_),
    .X(_03460_));
 sky130_fd_sc_hd__or2_2 _08540_ (.A(_02163_),
    .B(\rvsingle.dp.rf.rf[30][13] ),
    .X(_03461_));
 sky130_fd_sc_hd__o211a_2 _08541_ (.A1(_01440_),
    .A2(\rvsingle.dp.rf.rf[31][13] ),
    .B1(_02162_),
    .C1(_03461_),
    .X(_03462_));
 sky130_fd_sc_hd__or2_2 _08542_ (.A(_01349_),
    .B(\rvsingle.dp.rf.rf[28][13] ),
    .X(_03463_));
 sky130_fd_sc_hd__o211ai_2 _08543_ (.A1(\rvsingle.dp.rf.rf[29][13] ),
    .A2(_02275_),
    .B1(_01436_),
    .C1(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__nand2_2 _08544_ (.A(_03464_),
    .B(_02291_),
    .Y(_03465_));
 sky130_fd_sc_hd__o221ai_2 _08545_ (.A1(_01229_),
    .A2(_03460_),
    .B1(_03462_),
    .B2(_03465_),
    .C1(_02438_),
    .Y(_03466_));
 sky130_fd_sc_hd__o211ai_2 _08546_ (.A1(_03457_),
    .A2(_03459_),
    .B1(_03466_),
    .C1(_01187_),
    .Y(_03467_));
 sky130_fd_sc_hd__mux4_2 _08547_ (.A0(\rvsingle.dp.rf.rf[8][13] ),
    .A1(\rvsingle.dp.rf.rf[9][13] ),
    .A2(\rvsingle.dp.rf.rf[10][13] ),
    .A3(\rvsingle.dp.rf.rf[11][13] ),
    .S0(_01241_),
    .S1(_01953_),
    .X(_03468_));
 sky130_fd_sc_hd__mux2_2 _08548_ (.A0(\rvsingle.dp.rf.rf[12][13] ),
    .A1(\rvsingle.dp.rf.rf[13][13] ),
    .S(_01468_),
    .X(_03469_));
 sky130_fd_sc_hd__o21a_2 _08549_ (.A1(_01240_),
    .A2(\rvsingle.dp.rf.rf[14][13] ),
    .B1(_01454_),
    .X(_03470_));
 sky130_fd_sc_hd__o21a_2 _08550_ (.A1(_02929_),
    .A2(\rvsingle.dp.rf.rf[15][13] ),
    .B1(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__a211o_2 _08551_ (.A1(_03469_),
    .A2(_01716_),
    .B1(_01460_),
    .C1(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__o211ai_2 _08552_ (.A1(_01694_),
    .A2(_03468_),
    .B1(_01221_),
    .C1(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__mux4_2 _08553_ (.A0(\rvsingle.dp.rf.rf[0][13] ),
    .A1(\rvsingle.dp.rf.rf[1][13] ),
    .A2(\rvsingle.dp.rf.rf[2][13] ),
    .A3(\rvsingle.dp.rf.rf[3][13] ),
    .S0(_01241_),
    .S1(_01953_),
    .X(_03474_));
 sky130_fd_sc_hd__nor2_2 _08554_ (.A(_01463_),
    .B(\rvsingle.dp.rf.rf[6][13] ),
    .Y(_03475_));
 sky130_fd_sc_hd__o21ai_2 _08555_ (.A1(\rvsingle.dp.rf.rf[7][13] ),
    .A2(_02303_),
    .B1(_01199_),
    .Y(_03476_));
 sky130_fd_sc_hd__nor2_2 _08556_ (.A(_01463_),
    .B(\rvsingle.dp.rf.rf[4][13] ),
    .Y(_03477_));
 sky130_fd_sc_hd__o21ai_2 _08557_ (.A1(\rvsingle.dp.rf.rf[5][13] ),
    .A2(_01901_),
    .B1(_02285_),
    .Y(_03478_));
 sky130_fd_sc_hd__o221ai_2 _08558_ (.A1(_03475_),
    .A2(_03476_),
    .B1(_03477_),
    .B2(_03478_),
    .C1(_01702_),
    .Y(_03479_));
 sky130_fd_sc_hd__o211ai_2 _08559_ (.A1(_01694_),
    .A2(_03474_),
    .B1(_03479_),
    .C1(_01699_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand3_2 _08560_ (.A(_01316_),
    .B(_03473_),
    .C(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__o211ai_2 _08561_ (.A1(_01201_),
    .A2(_01351_),
    .B1(_03467_),
    .C1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__o21bai_2 _08562_ (.A1(_01184_),
    .A2(_03455_),
    .B1_N(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__mux2_2 _08563_ (.A0(\rvsingle.dp.rf.rf[0][12] ),
    .A1(\rvsingle.dp.rf.rf[1][12] ),
    .S(_01691_),
    .X(_03484_));
 sky130_fd_sc_hd__or2_2 _08564_ (.A(_01468_),
    .B(\rvsingle.dp.rf.rf[2][12] ),
    .X(_03485_));
 sky130_fd_sc_hd__o211a_2 _08565_ (.A1(_02303_),
    .A2(\rvsingle.dp.rf.rf[3][12] ),
    .B1(_01953_),
    .C1(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__a211oi_2 _08566_ (.A1(_03484_),
    .A2(_01309_),
    .B1(_01229_),
    .C1(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__mux4_2 _08567_ (.A0(\rvsingle.dp.rf.rf[4][12] ),
    .A1(\rvsingle.dp.rf.rf[5][12] ),
    .A2(\rvsingle.dp.rf.rf[6][12] ),
    .A3(\rvsingle.dp.rf.rf[7][12] ),
    .S0(_02450_),
    .S1(_01708_),
    .X(_03488_));
 sky130_fd_sc_hd__o21ai_2 _08568_ (.A1(_01207_),
    .A2(_03488_),
    .B1(_02447_),
    .Y(_03489_));
 sky130_fd_sc_hd__mux4_2 _08569_ (.A0(\rvsingle.dp.rf.rf[12][12] ),
    .A1(\rvsingle.dp.rf.rf[13][12] ),
    .A2(\rvsingle.dp.rf.rf[14][12] ),
    .A3(\rvsingle.dp.rf.rf[15][12] ),
    .S0(_02176_),
    .S1(_01696_),
    .X(_03490_));
 sky130_fd_sc_hd__nor2_2 _08570_ (.A(_01469_),
    .B(\rvsingle.dp.rf.rf[8][12] ),
    .Y(_03491_));
 sky130_fd_sc_hd__o21ai_2 _08571_ (.A1(\rvsingle.dp.rf.rf[9][12] ),
    .A2(_01295_),
    .B1(_02285_),
    .Y(_03492_));
 sky130_fd_sc_hd__o21a_2 _08572_ (.A1(_02450_),
    .A2(\rvsingle.dp.rf.rf[10][12] ),
    .B1(_01427_),
    .X(_03493_));
 sky130_fd_sc_hd__o21ai_2 _08573_ (.A1(\rvsingle.dp.rf.rf[11][12] ),
    .A2(_01901_),
    .B1(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__o211ai_2 _08574_ (.A1(_03491_),
    .A2(_03492_),
    .B1(_02543_),
    .C1(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__o211ai_2 _08575_ (.A1(_01422_),
    .A2(_03490_),
    .B1(_03495_),
    .C1(_01221_),
    .Y(_03496_));
 sky130_fd_sc_hd__o211a_2 _08576_ (.A1(_03487_),
    .A2(_03489_),
    .B1(_01315_),
    .C1(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__mux2_2 _08577_ (.A0(\rvsingle.dp.rf.rf[24][12] ),
    .A1(\rvsingle.dp.rf.rf[25][12] ),
    .S(_01691_),
    .X(_03498_));
 sky130_fd_sc_hd__or2_2 _08578_ (.A(_01462_),
    .B(\rvsingle.dp.rf.rf[26][12] ),
    .X(_03499_));
 sky130_fd_sc_hd__o211a_2 _08579_ (.A1(_02303_),
    .A2(\rvsingle.dp.rf.rf[27][12] ),
    .B1(_01199_),
    .C1(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__a211oi_2 _08580_ (.A1(_03498_),
    .A2(_01309_),
    .B1(_02302_),
    .C1(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__mux4_2 _08581_ (.A0(\rvsingle.dp.rf.rf[28][12] ),
    .A1(\rvsingle.dp.rf.rf[29][12] ),
    .A2(\rvsingle.dp.rf.rf[30][12] ),
    .A3(\rvsingle.dp.rf.rf[31][12] ),
    .S0(_01416_),
    .S1(_01300_),
    .X(_03502_));
 sky130_fd_sc_hd__o21ai_2 _08582_ (.A1(_01422_),
    .A2(_03502_),
    .B1(_01221_),
    .Y(_03503_));
 sky130_fd_sc_hd__mux4_2 _08583_ (.A0(\rvsingle.dp.rf.rf[16][12] ),
    .A1(\rvsingle.dp.rf.rf[17][12] ),
    .A2(\rvsingle.dp.rf.rf[18][12] ),
    .A3(\rvsingle.dp.rf.rf[19][12] ),
    .S0(_01730_),
    .S1(_01808_),
    .X(_03504_));
 sky130_fd_sc_hd__inv_2 _08584_ (.A(\rvsingle.dp.rf.rf[21][12] ),
    .Y(_03505_));
 sky130_fd_sc_hd__nor2_2 _08585_ (.A(_01328_),
    .B(\rvsingle.dp.rf.rf[20][12] ),
    .Y(_03506_));
 sky130_fd_sc_hd__a211o_2 _08586_ (.A1(_03505_),
    .A2(_01335_),
    .B1(_01727_),
    .C1(_03506_),
    .X(_03507_));
 sky130_fd_sc_hd__o21a_2 _08587_ (.A1(_01903_),
    .A2(\rvsingle.dp.rf.rf[22][12] ),
    .B1(_01243_),
    .X(_03508_));
 sky130_fd_sc_hd__o21ai_2 _08588_ (.A1(\rvsingle.dp.rf.rf[23][12] ),
    .A2(_01901_),
    .B1(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__a31oi_2 _08589_ (.A1(_03507_),
    .A2(_01702_),
    .A3(_03509_),
    .B1(_01446_),
    .Y(_03510_));
 sky130_fd_sc_hd__o21ai_2 _08590_ (.A1(_01694_),
    .A2(_03504_),
    .B1(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__o211ai_2 _08591_ (.A1(_03501_),
    .A2(_03503_),
    .B1(_02315_),
    .C1(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__nor3b_2 _08592_ (.A(_01452_),
    .B(_03497_),
    .C_N(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__o21bai_2 _08593_ (.A1(_02117_),
    .A2(\rvsingle.dp.rf.rf[8][12] ),
    .B1_N(_01530_),
    .Y(_03514_));
 sky130_fd_sc_hd__and2b_2 _08594_ (.A_N(\rvsingle.dp.rf.rf[9][12] ),
    .B(_03258_),
    .X(_03515_));
 sky130_fd_sc_hd__o21ai_2 _08595_ (.A1(_03514_),
    .A2(_03515_),
    .B1(_01131_),
    .Y(_03516_));
 sky130_fd_sc_hd__or2b_2 _08596_ (.A(\rvsingle.dp.rf.rf[11][12] ),
    .B_N(_01492_),
    .X(_03517_));
 sky130_fd_sc_hd__o211a_2 _08597_ (.A1(_01499_),
    .A2(\rvsingle.dp.rf.rf[10][12] ),
    .B1(_02059_),
    .C1(_03517_),
    .X(_03518_));
 sky130_fd_sc_hd__nor2_2 _08598_ (.A(_01630_),
    .B(\rvsingle.dp.rf.rf[12][12] ),
    .Y(_03519_));
 sky130_fd_sc_hd__and2b_2 _08599_ (.A_N(\rvsingle.dp.rf.rf[13][12] ),
    .B(_01618_),
    .X(_03520_));
 sky130_fd_sc_hd__or2b_2 _08600_ (.A(\rvsingle.dp.rf.rf[15][12] ),
    .B_N(_01566_),
    .X(_03521_));
 sky130_fd_sc_hd__o211ai_2 _08601_ (.A1(_01382_),
    .A2(\rvsingle.dp.rf.rf[14][12] ),
    .B1(_01777_),
    .C1(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__o311ai_2 _08602_ (.A1(_01620_),
    .A2(_03519_),
    .A3(_03520_),
    .B1(_02323_),
    .C1(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__o211ai_2 _08603_ (.A1(_03516_),
    .A2(_03518_),
    .B1(_01505_),
    .C1(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__inv_2 _08604_ (.A(\rvsingle.dp.rf.rf[5][12] ),
    .Y(_03525_));
 sky130_fd_sc_hd__nor2_2 _08605_ (.A(_01780_),
    .B(\rvsingle.dp.rf.rf[4][12] ),
    .Y(_03526_));
 sky130_fd_sc_hd__a211oi_2 _08606_ (.A1(_03525_),
    .A2(_01256_),
    .B1(_01531_),
    .C1(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__o21ai_2 _08607_ (.A1(_01558_),
    .A2(\rvsingle.dp.rf.rf[6][12] ),
    .B1(_01777_),
    .Y(_03528_));
 sky130_fd_sc_hd__and2b_2 _08608_ (.A_N(\rvsingle.dp.rf.rf[7][12] ),
    .B(_01650_),
    .X(_03529_));
 sky130_fd_sc_hd__o21ai_2 _08609_ (.A1(_03528_),
    .A2(_03529_),
    .B1(_02410_),
    .Y(_03530_));
 sky130_fd_sc_hd__nor2_2 _08610_ (.A(_01630_),
    .B(\rvsingle.dp.rf.rf[0][12] ),
    .Y(_03531_));
 sky130_fd_sc_hd__and2b_2 _08611_ (.A_N(\rvsingle.dp.rf.rf[1][12] ),
    .B(_01561_),
    .X(_03532_));
 sky130_fd_sc_hd__or2b_2 _08612_ (.A(\rvsingle.dp.rf.rf[3][12] ),
    .B_N(_01779_),
    .X(_03533_));
 sky130_fd_sc_hd__o211ai_2 _08613_ (.A1(_01382_),
    .A2(\rvsingle.dp.rf.rf[2][12] ),
    .B1(_01777_),
    .C1(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__o311ai_2 _08614_ (.A1(_01620_),
    .A2(_03531_),
    .A3(_03532_),
    .B1(_01131_),
    .C1(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__o211ai_2 _08615_ (.A1(_03527_),
    .A2(_03530_),
    .B1(_01156_),
    .C1(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand3_2 _08616_ (.A(_01377_),
    .B(_03524_),
    .C(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__nor2_2 _08617_ (.A(_01878_),
    .B(\rvsingle.dp.rf.rf[20][12] ),
    .Y(_03538_));
 sky130_fd_sc_hd__a211oi_2 _08618_ (.A1(_03505_),
    .A2(_01603_),
    .B1(_01660_),
    .C1(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__o21ai_2 _08619_ (.A1(_01382_),
    .A2(\rvsingle.dp.rf.rf[22][12] ),
    .B1(_02337_),
    .Y(_03540_));
 sky130_fd_sc_hd__and2b_2 _08620_ (.A_N(\rvsingle.dp.rf.rf[23][12] ),
    .B(_02005_),
    .X(_03541_));
 sky130_fd_sc_hd__o21ai_2 _08621_ (.A1(_03540_),
    .A2(_03541_),
    .B1(_01511_),
    .Y(_03542_));
 sky130_fd_sc_hd__nor2_2 _08622_ (.A(_01567_),
    .B(\rvsingle.dp.rf.rf[16][12] ),
    .Y(_03543_));
 sky130_fd_sc_hd__and2b_2 _08623_ (.A_N(\rvsingle.dp.rf.rf[17][12] ),
    .B(_03258_),
    .X(_03544_));
 sky130_fd_sc_hd__or2b_2 _08624_ (.A(\rvsingle.dp.rf.rf[19][12] ),
    .B_N(_02627_),
    .X(_03545_));
 sky130_fd_sc_hd__o211ai_2 _08625_ (.A1(_01545_),
    .A2(\rvsingle.dp.rf.rf[18][12] ),
    .B1(_02337_),
    .C1(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__o311ai_2 _08626_ (.A1(_01660_),
    .A2(_03543_),
    .A3(_03544_),
    .B1(_02351_),
    .C1(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__o211ai_2 _08627_ (.A1(_03539_),
    .A2(_03542_),
    .B1(_01156_),
    .C1(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__or2b_2 _08628_ (.A(\rvsingle.dp.rf.rf[29][12] ),
    .B_N(_01492_),
    .X(_03549_));
 sky130_fd_sc_hd__o211ai_2 _08629_ (.A1(_01137_),
    .A2(\rvsingle.dp.rf.rf[28][12] ),
    .B1(_03549_),
    .C1(_02485_),
    .Y(_03550_));
 sky130_fd_sc_hd__o21a_2 _08630_ (.A1(_01561_),
    .A2(\rvsingle.dp.rf.rf[30][12] ),
    .B1(_01530_),
    .X(_03551_));
 sky130_fd_sc_hd__o21ai_2 _08631_ (.A1(\rvsingle.dp.rf.rf[31][12] ),
    .A2(_01677_),
    .B1(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__nand3_2 _08632_ (.A(_03550_),
    .B(_02488_),
    .C(_03552_),
    .Y(_03553_));
 sky130_fd_sc_hd__and2b_2 _08633_ (.A_N(\rvsingle.dp.rf.rf[25][12] ),
    .B(_01769_),
    .X(_03554_));
 sky130_fd_sc_hd__o21ai_2 _08634_ (.A1(_01545_),
    .A2(\rvsingle.dp.rf.rf[24][12] ),
    .B1(_02395_),
    .Y(_03555_));
 sky130_fd_sc_hd__o21a_2 _08635_ (.A1(_01613_),
    .A2(\rvsingle.dp.rf.rf[26][12] ),
    .B1(_01551_),
    .X(_03556_));
 sky130_fd_sc_hd__o21ai_2 _08636_ (.A1(\rvsingle.dp.rf.rf[27][12] ),
    .A2(_01487_),
    .B1(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__o211ai_2 _08637_ (.A1(_03554_),
    .A2(_03555_),
    .B1(_02351_),
    .C1(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__nand3_2 _08638_ (.A(_03553_),
    .B(_03558_),
    .C(_02527_),
    .Y(_03559_));
 sky130_fd_sc_hd__nand3_2 _08639_ (.A(_03548_),
    .B(_01146_),
    .C(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__a31o_2 _08640_ (.A1(_02505_),
    .A2(_03537_),
    .A3(_03560_),
    .B1(_01177_),
    .X(_03561_));
 sky130_fd_sc_hd__o211ai_2 _08641_ (.A1(_01537_),
    .A2(_01171_),
    .B1(_01183_),
    .C1(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__a31oi_2 _08642_ (.A1(_02505_),
    .A2(_03537_),
    .A3(_03560_),
    .B1(_02375_),
    .Y(_03563_));
 sky130_fd_sc_hd__o22ai_2 _08643_ (.A1(_02473_),
    .A2(_02102_),
    .B1(_03142_),
    .B2(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand3_2 _08644_ (.A(_03513_),
    .B(_03562_),
    .C(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__o21ai_2 _08645_ (.A1(_01303_),
    .A2(_01351_),
    .B1(_03512_),
    .Y(_03566_));
 sky130_fd_sc_hd__o2bb2ai_2 _08646_ (.A1_N(_03562_),
    .A2_N(_03564_),
    .B1(_03497_),
    .B2(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__a31o_2 _08647_ (.A1(_01316_),
    .A2(_03473_),
    .A3(_03480_),
    .B1(_01452_),
    .X(_03568_));
 sky130_fd_sc_hd__inv_2 _08648_ (.A(_03467_),
    .Y(_03569_));
 sky130_fd_sc_hd__a31o_2 _08649_ (.A1(_02505_),
    .A2(_03452_),
    .A3(_03429_),
    .B1(_02375_),
    .X(_03570_));
 sky130_fd_sc_hd__a2bb2oi_2 _08650_ (.A1_N(_01960_),
    .A2_N(_02102_),
    .B1(_02261_),
    .B2(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__o22ai_2 _08651_ (.A1(_03568_),
    .A2(_03569_),
    .B1(_03454_),
    .B2(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__o2111ai_2 _08652_ (.A1(_03454_),
    .A2(_03483_),
    .B1(_03565_),
    .C1(_03567_),
    .D1(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__mux4_2 _08653_ (.A0(\rvsingle.dp.rf.rf[8][14] ),
    .A1(\rvsingle.dp.rf.rf[9][14] ),
    .A2(\rvsingle.dp.rf.rf[10][14] ),
    .A3(\rvsingle.dp.rf.rf[11][14] ),
    .S0(_01730_),
    .S1(_01953_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_2 _08654_ (.A0(\rvsingle.dp.rf.rf[12][14] ),
    .A1(\rvsingle.dp.rf.rf[13][14] ),
    .S(_01828_),
    .X(_03575_));
 sky130_fd_sc_hd__or2_2 _08655_ (.A(_01425_),
    .B(\rvsingle.dp.rf.rf[14][14] ),
    .X(_03576_));
 sky130_fd_sc_hd__o211a_2 _08656_ (.A1(_01423_),
    .A2(\rvsingle.dp.rf.rf[15][14] ),
    .B1(_01427_),
    .C1(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__a211o_2 _08657_ (.A1(_03575_),
    .A2(_01716_),
    .B1(_01460_),
    .C1(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__o211ai_2 _08658_ (.A1(_01694_),
    .A2(_03574_),
    .B1(_03578_),
    .C1(_01221_),
    .Y(_03579_));
 sky130_fd_sc_hd__mux4_2 _08659_ (.A0(\rvsingle.dp.rf.rf[0][14] ),
    .A1(\rvsingle.dp.rf.rf[1][14] ),
    .A2(\rvsingle.dp.rf.rf[2][14] ),
    .A3(\rvsingle.dp.rf.rf[3][14] ),
    .S0(_01730_),
    .S1(_01433_),
    .X(_03580_));
 sky130_fd_sc_hd__mux2_2 _08660_ (.A0(\rvsingle.dp.rf.rf[4][14] ),
    .A1(\rvsingle.dp.rf.rf[5][14] ),
    .S(_01468_),
    .X(_03581_));
 sky130_fd_sc_hd__or2_2 _08661_ (.A(_01425_),
    .B(\rvsingle.dp.rf.rf[6][14] ),
    .X(_03582_));
 sky130_fd_sc_hd__o211a_2 _08662_ (.A1(_02929_),
    .A2(\rvsingle.dp.rf.rf[7][14] ),
    .B1(_01427_),
    .C1(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__a211o_2 _08663_ (.A1(_03581_),
    .A2(_01716_),
    .B1(_01460_),
    .C1(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__o211ai_2 _08664_ (.A1(_03580_),
    .A2(_01445_),
    .B1(_01699_),
    .C1(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__nand3_2 _08665_ (.A(_01316_),
    .B(_03579_),
    .C(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__mux4_2 _08666_ (.A0(\rvsingle.dp.rf.rf[20][14] ),
    .A1(\rvsingle.dp.rf.rf[21][14] ),
    .A2(\rvsingle.dp.rf.rf[22][14] ),
    .A3(\rvsingle.dp.rf.rf[23][14] ),
    .S0(_01241_),
    .S1(_01953_),
    .X(_03587_));
 sky130_fd_sc_hd__nor2_2 _08667_ (.A(_02093_),
    .B(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__mux4_2 _08668_ (.A0(\rvsingle.dp.rf.rf[16][14] ),
    .A1(\rvsingle.dp.rf.rf[17][14] ),
    .A2(\rvsingle.dp.rf.rf[18][14] ),
    .A3(\rvsingle.dp.rf.rf[19][14] ),
    .S0(_01426_),
    .S1(_02162_),
    .X(_03589_));
 sky130_fd_sc_hd__o21ai_2 _08669_ (.A1(_01711_),
    .A2(_03589_),
    .B1(_01699_),
    .Y(_03590_));
 sky130_fd_sc_hd__mux4_2 _08670_ (.A0(\rvsingle.dp.rf.rf[24][14] ),
    .A1(\rvsingle.dp.rf.rf[25][14] ),
    .A2(\rvsingle.dp.rf.rf[26][14] ),
    .A3(\rvsingle.dp.rf.rf[27][14] ),
    .S0(_01426_),
    .S1(_01433_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_2 _08671_ (.A0(\rvsingle.dp.rf.rf[28][14] ),
    .A1(\rvsingle.dp.rf.rf[29][14] ),
    .S(_01191_),
    .X(_03592_));
 sky130_fd_sc_hd__or2b_2 _08672_ (.A(\rvsingle.dp.rf.rf[31][14] ),
    .B_N(_01425_),
    .X(_03593_));
 sky130_fd_sc_hd__o211a_2 _08673_ (.A1(_02450_),
    .A2(\rvsingle.dp.rf.rf[30][14] ),
    .B1(_01427_),
    .C1(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__a211o_2 _08674_ (.A1(_03592_),
    .A2(_01716_),
    .B1(_01460_),
    .C1(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__o211ai_2 _08675_ (.A1(_01711_),
    .A2(_03591_),
    .B1(_03595_),
    .C1(_01221_),
    .Y(_03596_));
 sky130_fd_sc_hd__o211ai_2 _08676_ (.A1(_03588_),
    .A2(_03590_),
    .B1(_02315_),
    .C1(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__nor2_2 _08677_ (.A(_01619_),
    .B(\rvsingle.dp.rf.rf[30][14] ),
    .Y(_03598_));
 sky130_fd_sc_hd__o21ai_2 _08678_ (.A1(\rvsingle.dp.rf.rf[31][14] ),
    .A2(_01677_),
    .B1(_02320_),
    .Y(_03599_));
 sky130_fd_sc_hd__or2_2 _08679_ (.A(_01267_),
    .B(\rvsingle.dp.rf.rf[28][14] ),
    .X(_03600_));
 sky130_fd_sc_hd__o211ai_2 _08680_ (.A1(\rvsingle.dp.rf.rf[29][14] ),
    .A2(_02481_),
    .B1(_01496_),
    .C1(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__o211ai_2 _08681_ (.A1(_03598_),
    .A2(_03599_),
    .B1(_03601_),
    .C1(_01617_),
    .Y(_03602_));
 sky130_fd_sc_hd__nor2_2 _08682_ (.A(_01780_),
    .B(\rvsingle.dp.rf.rf[24][14] ),
    .Y(_03603_));
 sky130_fd_sc_hd__and2b_2 _08683_ (.A_N(\rvsingle.dp.rf.rf[25][14] ),
    .B(_01769_),
    .X(_03604_));
 sky130_fd_sc_hd__o21a_2 _08684_ (.A1(_01613_),
    .A2(\rvsingle.dp.rf.rf[26][14] ),
    .B1(_01551_),
    .X(_03605_));
 sky130_fd_sc_hd__o21ai_2 _08685_ (.A1(\rvsingle.dp.rf.rf[27][14] ),
    .A2(_01487_),
    .B1(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__o311ai_2 _08686_ (.A1(_01605_),
    .A2(_03603_),
    .A3(_03604_),
    .B1(_02351_),
    .C1(_03606_),
    .Y(_03607_));
 sky130_fd_sc_hd__nand3_2 _08687_ (.A(_03602_),
    .B(_03607_),
    .C(_02527_),
    .Y(_03608_));
 sky130_fd_sc_hd__nor2_2 _08688_ (.A(_01382_),
    .B(\rvsingle.dp.rf.rf[16][14] ),
    .Y(_03609_));
 sky130_fd_sc_hd__and2b_2 _08689_ (.A_N(\rvsingle.dp.rf.rf[17][14] ),
    .B(_01255_),
    .X(_03610_));
 sky130_fd_sc_hd__or2b_2 _08690_ (.A(\rvsingle.dp.rf.rf[19][14] ),
    .B_N(_01779_),
    .X(_03611_));
 sky130_fd_sc_hd__o211ai_2 _08691_ (.A1(_01567_),
    .A2(\rvsingle.dp.rf.rf[18][14] ),
    .B1(_02031_),
    .C1(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__o311ai_2 _08692_ (.A1(_01531_),
    .A2(_03609_),
    .A3(_03610_),
    .B1(_01131_),
    .C1(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__nor2_2 _08693_ (.A(_01763_),
    .B(\rvsingle.dp.rf.rf[22][14] ),
    .Y(_03614_));
 sky130_fd_sc_hd__and2b_2 _08694_ (.A_N(\rvsingle.dp.rf.rf[23][14] ),
    .B(_03258_),
    .X(_03615_));
 sky130_fd_sc_hd__o21ba_2 _08695_ (.A1(_01267_),
    .A2(\rvsingle.dp.rf.rf[20][14] ),
    .B1_N(_01258_),
    .X(_03616_));
 sky130_fd_sc_hd__o21ai_2 _08696_ (.A1(_01539_),
    .A2(\rvsingle.dp.rf.rf[21][14] ),
    .B1(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__o311ai_2 _08697_ (.A1(_02485_),
    .A2(_03614_),
    .A3(_03615_),
    .B1(_02410_),
    .C1(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand3_2 _08698_ (.A(_01853_),
    .B(_03613_),
    .C(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__nand3_2 _08699_ (.A(_03608_),
    .B(_03619_),
    .C(_01146_),
    .Y(_03620_));
 sky130_fd_sc_hd__nor2_2 _08700_ (.A(_01137_),
    .B(\rvsingle.dp.rf.rf[10][14] ),
    .Y(_03621_));
 sky130_fd_sc_hd__o21ai_2 _08701_ (.A1(\rvsingle.dp.rf.rf[11][14] ),
    .A2(_01487_),
    .B1(_01523_),
    .Y(_03622_));
 sky130_fd_sc_hd__or2b_2 _08702_ (.A(\rvsingle.dp.rf.rf[9][14] ),
    .B_N(_01498_),
    .X(_03623_));
 sky130_fd_sc_hd__o211ai_2 _08703_ (.A1(_01499_),
    .A2(\rvsingle.dp.rf.rf[8][14] ),
    .B1(_03623_),
    .C1(_01496_),
    .Y(_03624_));
 sky130_fd_sc_hd__o211ai_2 _08704_ (.A1(_03621_),
    .A2(_03622_),
    .B1(_03624_),
    .C1(_02483_),
    .Y(_03625_));
 sky130_fd_sc_hd__o21ba_2 _08705_ (.A1(_01255_),
    .A2(\rvsingle.dp.rf.rf[12][14] ),
    .B1_N(_01551_),
    .X(_03626_));
 sky130_fd_sc_hd__o21ai_2 _08706_ (.A1(_01677_),
    .A2(\rvsingle.dp.rf.rf[13][14] ),
    .B1(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__o21a_2 _08707_ (.A1(_01618_),
    .A2(\rvsingle.dp.rf.rf[14][14] ),
    .B1(_01530_),
    .X(_03628_));
 sky130_fd_sc_hd__o21ai_2 _08708_ (.A1(\rvsingle.dp.rf.rf[15][14] ),
    .A2(_02481_),
    .B1(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__nand3_2 _08709_ (.A(_03627_),
    .B(_02488_),
    .C(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__nand3_2 _08710_ (.A(_03625_),
    .B(_02527_),
    .C(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__nor2_2 _08711_ (.A(_01567_),
    .B(\rvsingle.dp.rf.rf[0][14] ),
    .Y(_03632_));
 sky130_fd_sc_hd__and2b_2 _08712_ (.A_N(\rvsingle.dp.rf.rf[1][14] ),
    .B(_03258_),
    .X(_03633_));
 sky130_fd_sc_hd__or2b_2 _08713_ (.A(\rvsingle.dp.rf.rf[3][14] ),
    .B_N(_01877_),
    .X(_03634_));
 sky130_fd_sc_hd__o211ai_2 _08714_ (.A1(_01545_),
    .A2(\rvsingle.dp.rf.rf[2][14] ),
    .B1(_02337_),
    .C1(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__o311ai_2 _08715_ (.A1(_01531_),
    .A2(_03632_),
    .A3(_03633_),
    .B1(_02351_),
    .C1(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__nor2_2 _08716_ (.A(_01567_),
    .B(\rvsingle.dp.rf.rf[4][14] ),
    .Y(_03637_));
 sky130_fd_sc_hd__and2b_2 _08717_ (.A_N(\rvsingle.dp.rf.rf[5][14] ),
    .B(_03258_),
    .X(_03638_));
 sky130_fd_sc_hd__or2b_2 _08718_ (.A(\rvsingle.dp.rf.rf[7][14] ),
    .B_N(_01877_),
    .X(_03639_));
 sky130_fd_sc_hd__o211ai_2 _08719_ (.A1(_01545_),
    .A2(\rvsingle.dp.rf.rf[6][14] ),
    .B1(_02337_),
    .C1(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__o311ai_2 _08720_ (.A1(_01660_),
    .A2(_03637_),
    .A3(_03638_),
    .B1(_02410_),
    .C1(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__nand3_2 _08721_ (.A(_01853_),
    .B(_03636_),
    .C(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__nand3_2 _08722_ (.A(_01377_),
    .B(_03631_),
    .C(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__o211ai_2 _08723_ (.A1(_01962_),
    .A2(_01128_),
    .B1(_03620_),
    .C1(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__o221ai_2 _08724_ (.A1(_02473_),
    .A2(_02318_),
    .B1(_01961_),
    .B2(_03644_),
    .C1(_01580_),
    .Y(_03645_));
 sky130_fd_sc_hd__a31o_2 _08725_ (.A1(_02505_),
    .A2(_03643_),
    .A3(_03620_),
    .B1(_02375_),
    .X(_03646_));
 sky130_fd_sc_hd__nand3_2 _08726_ (.A(_03646_),
    .B(_01183_),
    .C(_02261_),
    .Y(_03647_));
 sky130_fd_sc_hd__a32o_2 _08727_ (.A1(_01248_),
    .A2(_03586_),
    .A3(_03597_),
    .B1(_03645_),
    .B2(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__o311a_2 _08728_ (.A1(_01338_),
    .A2(_01245_),
    .A3(_01201_),
    .B1(_03597_),
    .C1(_03586_),
    .X(_03649_));
 sky130_fd_sc_hd__nand3_2 _08729_ (.A(_03647_),
    .B(_03649_),
    .C(_03645_),
    .Y(_03650_));
 sky130_fd_sc_hd__nor2_2 _08730_ (.A(_01595_),
    .B(\rvsingle.dp.rf.rf[18][15] ),
    .Y(_03651_));
 sky130_fd_sc_hd__o21ai_2 _08731_ (.A1(\rvsingle.dp.rf.rf[19][15] ),
    .A2(_02478_),
    .B1(_01490_),
    .Y(_03652_));
 sky130_fd_sc_hd__or2b_2 _08732_ (.A(\rvsingle.dp.rf.rf[17][15] ),
    .B_N(_01877_),
    .X(_03653_));
 sky130_fd_sc_hd__o211ai_2 _08733_ (.A1(_01878_),
    .A2(\rvsingle.dp.rf.rf[16][15] ),
    .B1(_03653_),
    .C1(_02395_),
    .Y(_03654_));
 sky130_fd_sc_hd__o211ai_2 _08734_ (.A1(_03651_),
    .A2(_03652_),
    .B1(_03654_),
    .C1(_02483_),
    .Y(_03655_));
 sky130_fd_sc_hd__nor2_2 _08735_ (.A(_01595_),
    .B(\rvsingle.dp.rf.rf[22][15] ),
    .Y(_03656_));
 sky130_fd_sc_hd__o21ai_2 _08736_ (.A1(\rvsingle.dp.rf.rf[23][15] ),
    .A2(_02478_),
    .B1(_01490_),
    .Y(_03657_));
 sky130_fd_sc_hd__or2b_2 _08737_ (.A(\rvsingle.dp.rf.rf[21][15] ),
    .B_N(_01877_),
    .X(_03658_));
 sky130_fd_sc_hd__o211ai_2 _08738_ (.A1(_01878_),
    .A2(\rvsingle.dp.rf.rf[20][15] ),
    .B1(_03658_),
    .C1(_02395_),
    .Y(_03659_));
 sky130_fd_sc_hd__o211ai_2 _08739_ (.A1(_03656_),
    .A2(_03657_),
    .B1(_03659_),
    .C1(_02488_),
    .Y(_03660_));
 sky130_fd_sc_hd__nand3_2 _08740_ (.A(_01853_),
    .B(_03655_),
    .C(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__nor2_2 _08741_ (.A(_01137_),
    .B(\rvsingle.dp.rf.rf[30][15] ),
    .Y(_03662_));
 sky130_fd_sc_hd__o21ai_2 _08742_ (.A1(\rvsingle.dp.rf.rf[31][15] ),
    .A2(_01487_),
    .B1(_01523_),
    .Y(_03663_));
 sky130_fd_sc_hd__or2b_2 _08743_ (.A(\rvsingle.dp.rf.rf[29][15] ),
    .B_N(_02627_),
    .X(_03664_));
 sky130_fd_sc_hd__o211ai_2 _08744_ (.A1(_01499_),
    .A2(\rvsingle.dp.rf.rf[28][15] ),
    .B1(_03664_),
    .C1(_01496_),
    .Y(_03665_));
 sky130_fd_sc_hd__o211ai_2 _08745_ (.A1(_03662_),
    .A2(_03663_),
    .B1(_03665_),
    .C1(_02488_),
    .Y(_03666_));
 sky130_fd_sc_hd__nor2_2 _08746_ (.A(_01382_),
    .B(\rvsingle.dp.rf.rf[24][15] ),
    .Y(_03667_));
 sky130_fd_sc_hd__and2b_2 _08747_ (.A_N(\rvsingle.dp.rf.rf[25][15] ),
    .B(_01255_),
    .X(_03668_));
 sky130_fd_sc_hd__o21a_2 _08748_ (.A1(_01594_),
    .A2(\rvsingle.dp.rf.rf[26][15] ),
    .B1(_01489_),
    .X(_03669_));
 sky130_fd_sc_hd__o21ai_2 _08749_ (.A1(\rvsingle.dp.rf.rf[27][15] ),
    .A2(_01508_),
    .B1(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__o311ai_2 _08750_ (.A1(_01531_),
    .A2(_03667_),
    .A3(_03668_),
    .B1(_01131_),
    .C1(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__nand3_2 _08751_ (.A(_03666_),
    .B(_03671_),
    .C(_02527_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand3_2 _08752_ (.A(_03661_),
    .B(_01146_),
    .C(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__or2b_2 _08753_ (.A(\rvsingle.dp.rf.rf[11][15] ),
    .B_N(_01136_),
    .X(_03674_));
 sky130_fd_sc_hd__o211a_2 _08754_ (.A1(_01513_),
    .A2(\rvsingle.dp.rf.rf[10][15] ),
    .B1(_02059_),
    .C1(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__o21ba_2 _08755_ (.A1(_01561_),
    .A2(\rvsingle.dp.rf.rf[8][15] ),
    .B1_N(_01489_),
    .X(_03676_));
 sky130_fd_sc_hd__or2b_2 _08756_ (.A(\rvsingle.dp.rf.rf[9][15] ),
    .B_N(_01613_),
    .X(_03677_));
 sky130_fd_sc_hd__a21o_2 _08757_ (.A1(_03676_),
    .A2(_03677_),
    .B1(_01111_),
    .X(_03678_));
 sky130_fd_sc_hd__nor2_2 _08758_ (.A(_01513_),
    .B(\rvsingle.dp.rf.rf[14][15] ),
    .Y(_03679_));
 sky130_fd_sc_hd__o21ai_2 _08759_ (.A1(\rvsingle.dp.rf.rf[15][15] ),
    .A2(_01508_),
    .B1(_02059_),
    .Y(_03680_));
 sky130_fd_sc_hd__or2_2 _08760_ (.A(_01498_),
    .B(\rvsingle.dp.rf.rf[12][15] ),
    .X(_03681_));
 sky130_fd_sc_hd__o211ai_2 _08761_ (.A1(\rvsingle.dp.rf.rf[13][15] ),
    .A2(_01487_),
    .B1(_02395_),
    .C1(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__o211ai_2 _08762_ (.A1(_03679_),
    .A2(_03680_),
    .B1(_01511_),
    .C1(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__o211ai_2 _08763_ (.A1(_03675_),
    .A2(_03678_),
    .B1(_02527_),
    .C1(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__nor2_2 _08764_ (.A(_01595_),
    .B(\rvsingle.dp.rf.rf[0][15] ),
    .Y(_03685_));
 sky130_fd_sc_hd__o21bai_2 _08765_ (.A1(\rvsingle.dp.rf.rf[1][15] ),
    .A2(_02478_),
    .B1_N(_01647_),
    .Y(_03686_));
 sky130_fd_sc_hd__or2_2 _08766_ (.A(_01498_),
    .B(\rvsingle.dp.rf.rf[2][15] ),
    .X(_03687_));
 sky130_fd_sc_hd__o211ai_2 _08767_ (.A1(_02478_),
    .A2(\rvsingle.dp.rf.rf[3][15] ),
    .B1(_01490_),
    .C1(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__o211ai_2 _08768_ (.A1(_03685_),
    .A2(_03686_),
    .B1(_02351_),
    .C1(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__nor2_2 _08769_ (.A(_01545_),
    .B(\rvsingle.dp.rf.rf[4][15] ),
    .Y(_03690_));
 sky130_fd_sc_hd__and2b_2 _08770_ (.A_N(\rvsingle.dp.rf.rf[5][15] ),
    .B(_01602_),
    .X(_03691_));
 sky130_fd_sc_hd__or2b_2 _08771_ (.A(\rvsingle.dp.rf.rf[7][15] ),
    .B_N(_02627_),
    .X(_03692_));
 sky130_fd_sc_hd__o211ai_2 _08772_ (.A1(_02030_),
    .A2(\rvsingle.dp.rf.rf[6][15] ),
    .B1(_02337_),
    .C1(_03692_),
    .Y(_03693_));
 sky130_fd_sc_hd__o311ai_2 _08773_ (.A1(_01660_),
    .A2(_03690_),
    .A3(_03691_),
    .B1(_02410_),
    .C1(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__nand3_2 _08774_ (.A(_01853_),
    .B(_03689_),
    .C(_03694_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand3_2 _08775_ (.A(_01593_),
    .B(_03684_),
    .C(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__o211ai_2 _08776_ (.A1(_01962_),
    .A2(_01128_),
    .B1(_03673_),
    .C1(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__nand2_2 _08777_ (.A(_03697_),
    .B(_01537_),
    .Y(_03698_));
 sky130_fd_sc_hd__o211ai_2 _08778_ (.A1(_01084_),
    .A2(_01171_),
    .B1(_01584_),
    .C1(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__mux4_2 _08779_ (.A0(\rvsingle.dp.rf.rf[24][15] ),
    .A1(\rvsingle.dp.rf.rf[25][15] ),
    .A2(\rvsingle.dp.rf.rf[26][15] ),
    .A3(\rvsingle.dp.rf.rf[27][15] ),
    .S0(_01691_),
    .S1(_01244_),
    .X(_03700_));
 sky130_fd_sc_hd__mux2_2 _08780_ (.A0(\rvsingle.dp.rf.rf[30][15] ),
    .A1(\rvsingle.dp.rf.rf[31][15] ),
    .S(_01903_),
    .X(_03701_));
 sky130_fd_sc_hd__or2_2 _08781_ (.A(_01240_),
    .B(\rvsingle.dp.rf.rf[28][15] ),
    .X(_03702_));
 sky130_fd_sc_hd__o211a_2 _08782_ (.A1(\rvsingle.dp.rf.rf[29][15] ),
    .A2(_02929_),
    .B1(_01307_),
    .C1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__a211o_2 _08783_ (.A1(_01471_),
    .A2(_03701_),
    .B1(_02543_),
    .C1(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__o211ai_2 _08784_ (.A1(_01445_),
    .A2(_03700_),
    .B1(_01447_),
    .C1(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__mux4_2 _08785_ (.A0(\rvsingle.dp.rf.rf[20][15] ),
    .A1(\rvsingle.dp.rf.rf[21][15] ),
    .A2(\rvsingle.dp.rf.rf[22][15] ),
    .A3(\rvsingle.dp.rf.rf[23][15] ),
    .S0(_01691_),
    .S1(_01244_),
    .X(_03706_));
 sky130_fd_sc_hd__or2_2 _08786_ (.A(_02440_),
    .B(\rvsingle.dp.rf.rf[16][15] ),
    .X(_03707_));
 sky130_fd_sc_hd__o211ai_2 _08787_ (.A1(\rvsingle.dp.rf.rf[17][15] ),
    .A2(_01424_),
    .B1(_02285_),
    .C1(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__o21a_2 _08788_ (.A1(_01426_),
    .A2(\rvsingle.dp.rf.rf[18][15] ),
    .B1(_01427_),
    .X(_03709_));
 sky130_fd_sc_hd__o21ai_2 _08789_ (.A1(\rvsingle.dp.rf.rf[19][15] ),
    .A2(_01424_),
    .B1(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__a31oi_2 _08790_ (.A1(_01721_),
    .A2(_03708_),
    .A3(_03710_),
    .B1(_01446_),
    .Y(_03711_));
 sky130_fd_sc_hd__o21ai_2 _08791_ (.A1(_01461_),
    .A2(_03706_),
    .B1(_03711_),
    .Y(_03712_));
 sky130_fd_sc_hd__nand3_2 _08792_ (.A(_03705_),
    .B(_03712_),
    .C(_02315_),
    .Y(_03713_));
 sky130_fd_sc_hd__mux4_2 _08793_ (.A0(\rvsingle.dp.rf.rf[12][15] ),
    .A1(\rvsingle.dp.rf.rf[13][15] ),
    .A2(\rvsingle.dp.rf.rf[14][15] ),
    .A3(\rvsingle.dp.rf.rf[15][15] ),
    .S0(_01335_),
    .S1(_01199_),
    .X(_03714_));
 sky130_fd_sc_hd__mux2_2 _08794_ (.A0(\rvsingle.dp.rf.rf[8][15] ),
    .A1(\rvsingle.dp.rf.rf[9][15] ),
    .S(_02440_),
    .X(_03715_));
 sky130_fd_sc_hd__or2_2 _08795_ (.A(_01240_),
    .B(\rvsingle.dp.rf.rf[10][15] ),
    .X(_03716_));
 sky130_fd_sc_hd__o211a_2 _08796_ (.A1(_02929_),
    .A2(\rvsingle.dp.rf.rf[11][15] ),
    .B1(_01727_),
    .C1(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__a211o_2 _08797_ (.A1(_03715_),
    .A2(_01689_),
    .B1(_02273_),
    .C1(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__o211ai_2 _08798_ (.A1(_01461_),
    .A2(_03714_),
    .B1(_03718_),
    .C1(_01447_),
    .Y(_03719_));
 sky130_fd_sc_hd__mux4_2 _08799_ (.A0(\rvsingle.dp.rf.rf[4][15] ),
    .A1(\rvsingle.dp.rf.rf[5][15] ),
    .A2(\rvsingle.dp.rf.rf[6][15] ),
    .A3(\rvsingle.dp.rf.rf[7][15] ),
    .S0(_01335_),
    .S1(_01244_),
    .X(_03720_));
 sky130_fd_sc_hd__mux2_2 _08800_ (.A0(\rvsingle.dp.rf.rf[0][15] ),
    .A1(\rvsingle.dp.rf.rf[1][15] ),
    .S(_02440_),
    .X(_03721_));
 sky130_fd_sc_hd__or2_2 _08801_ (.A(_01240_),
    .B(\rvsingle.dp.rf.rf[2][15] ),
    .X(_03722_));
 sky130_fd_sc_hd__o211a_2 _08802_ (.A1(_02929_),
    .A2(\rvsingle.dp.rf.rf[3][15] ),
    .B1(_01727_),
    .C1(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__a211o_2 _08803_ (.A1(_03721_),
    .A2(_01689_),
    .B1(_02273_),
    .C1(_03723_),
    .X(_03724_));
 sky130_fd_sc_hd__o211ai_2 _08804_ (.A1(_01461_),
    .A2(_03720_),
    .B1(_03724_),
    .C1(_01218_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand3_2 _08805_ (.A(_01316_),
    .B(_03719_),
    .C(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__o311a_2 _08806_ (.A1(_01338_),
    .A2(_01201_),
    .A3(_01245_),
    .B1(_03713_),
    .C1(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__o221ai_2 _08807_ (.A1(_01960_),
    .A2(_02102_),
    .B1(_01961_),
    .B2(_03697_),
    .C1(_01580_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand3_2 _08808_ (.A(_03699_),
    .B(_03727_),
    .C(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand4_2 _08809_ (.A(_03696_),
    .B(_01481_),
    .C(_02505_),
    .D(_03673_),
    .Y(_03730_));
 sky130_fd_sc_hd__o211a_2 _08810_ (.A1(_02473_),
    .A2(_02318_),
    .B1(_01580_),
    .C1(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__a21oi_2 _08811_ (.A1(_01587_),
    .A2(_03730_),
    .B1(_01486_),
    .Y(_03732_));
 sky130_fd_sc_hd__o211ai_2 _08812_ (.A1(_01202_),
    .A2(_01351_),
    .B1(_03713_),
    .C1(_03726_),
    .Y(_03733_));
 sky130_fd_sc_hd__o21ai_2 _08813_ (.A1(_03731_),
    .A2(_03732_),
    .B1(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand4_2 _08814_ (.A(_03648_),
    .B(_03650_),
    .C(_03729_),
    .D(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__nor4_2 _08815_ (.A(_03231_),
    .B(_03406_),
    .C(_03573_),
    .D(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__o2111a_2 _08816_ (.A1(_03454_),
    .A2(_03483_),
    .B1(_03565_),
    .C1(_03567_),
    .D1(_03572_),
    .X(_03737_));
 sky130_fd_sc_hd__a21oi_2 _08817_ (.A1(_03645_),
    .A2(_03647_),
    .B1(_03649_),
    .Y(_03738_));
 sky130_fd_sc_hd__and3_2 _08818_ (.A(_03647_),
    .B(_03649_),
    .C(_03645_),
    .X(_03739_));
 sky130_fd_sc_hd__nor2_2 _08819_ (.A(_03738_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__a21oi_2 _08820_ (.A1(_03697_),
    .A2(_01085_),
    .B1(_01837_),
    .Y(_03741_));
 sky130_fd_sc_hd__a211oi_2 _08821_ (.A1(_03741_),
    .A2(_02261_),
    .B1(_03733_),
    .C1(_03731_),
    .Y(_03742_));
 sky130_fd_sc_hd__a21oi_2 _08822_ (.A1(_03728_),
    .A2(_03699_),
    .B1(_03727_),
    .Y(_03743_));
 sky130_fd_sc_hd__nor2_2 _08823_ (.A(_03742_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand3_2 _08824_ (.A(_03737_),
    .B(_03740_),
    .C(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__o211a_2 _08825_ (.A1(_03143_),
    .A2(_03141_),
    .B1(_03227_),
    .C1(_03221_),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_2 _08826_ (.A(_03397_),
    .B(_03382_),
    .Y(_03747_));
 sky130_fd_sc_hd__a2bb2oi_2 _08827_ (.A1_N(_02469_),
    .A2_N(_03747_),
    .B1(_03404_),
    .B2(_03402_),
    .Y(_03748_));
 sky130_fd_sc_hd__a21oi_2 _08828_ (.A1(_03313_),
    .A2(_03405_),
    .B1(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__a31o_2 _08829_ (.A1(_01153_),
    .A2(_03110_),
    .A3(_03087_),
    .B1(_01178_),
    .X(_03750_));
 sky130_fd_sc_hd__o211ai_2 _08830_ (.A1(_01482_),
    .A2(_01171_),
    .B1(_01584_),
    .C1(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__a2bb2oi_2 _08831_ (.A1_N(_02469_),
    .A2_N(_03228_),
    .B1(_03112_),
    .B2(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__o22ai_2 _08832_ (.A1(_03143_),
    .A2(_03141_),
    .B1(_03227_),
    .B2(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__a31oi_2 _08833_ (.A1(_03746_),
    .A2(_03749_),
    .A3(_03230_),
    .B1(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__o21ai_2 _08834_ (.A1(_03454_),
    .A2(_03483_),
    .B1(_03565_),
    .Y(_03755_));
 sky130_fd_sc_hd__o21ai_2 _08835_ (.A1(_03650_),
    .A2(_03743_),
    .B1(_03729_),
    .Y(_03756_));
 sky130_fd_sc_hd__a41oi_2 _08836_ (.A1(_03740_),
    .A2(_03744_),
    .A3(_03755_),
    .A4(_03572_),
    .B1(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__o21ai_2 _08837_ (.A1(_03745_),
    .A2(_03754_),
    .B1(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__a21oi_2 _08838_ (.A1(_03064_),
    .A2(_03736_),
    .B1(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__nand4_2 _08839_ (.A(_02015_),
    .B(_02016_),
    .C(_02098_),
    .D(_02100_),
    .Y(_03760_));
 sky130_fd_sc_hd__a21o_2 _08840_ (.A1(_02150_),
    .A2(_01482_),
    .B1(_01486_),
    .X(_03761_));
 sky130_fd_sc_hd__o21a_2 _08841_ (.A1(_03142_),
    .A2(_03761_),
    .B1(_02151_),
    .X(_03762_));
 sky130_fd_sc_hd__a21oi_2 _08842_ (.A1(_01581_),
    .A2(_02262_),
    .B1(_01837_),
    .Y(_03763_));
 sky130_fd_sc_hd__o31ai_2 _08843_ (.A1(_02211_),
    .A2(_02263_),
    .A3(_03763_),
    .B1(_02183_),
    .Y(_03764_));
 sky130_fd_sc_hd__o21ai_2 _08844_ (.A1(_02181_),
    .A2(_03762_),
    .B1(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__a21oi_2 _08845_ (.A1(_02012_),
    .A2(_02014_),
    .B1(_01959_),
    .Y(_03766_));
 sky130_fd_sc_hd__o21a_2 _08846_ (.A1(_03766_),
    .A2(_02100_),
    .B1(_02015_),
    .X(_03767_));
 sky130_fd_sc_hd__o21ai_2 _08847_ (.A1(_03760_),
    .A2(_03765_),
    .B1(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__nand2_2 _08848_ (.A(_01931_),
    .B(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__o22a_2 _08849_ (.A1(_01453_),
    .A2(_01480_),
    .B1(_01579_),
    .B2(_01582_),
    .X(_03770_));
 sky130_fd_sc_hd__a2111o_2 _08850_ (.A1(_01589_),
    .A2(_01739_),
    .B1(_03770_),
    .C1(_01840_),
    .D1(_01930_),
    .X(_03771_));
 sky130_fd_sc_hd__o21ba_2 _08851_ (.A1(_01838_),
    .A2(_01804_),
    .B1_N(_01834_),
    .X(_03772_));
 sky130_fd_sc_hd__o21a_2 _08852_ (.A1(_01927_),
    .A2(_03772_),
    .B1(_01836_),
    .X(_03773_));
 sky130_fd_sc_hd__nand3_2 _08853_ (.A(_03769_),
    .B(_03771_),
    .C(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__o21bai_2 _08854_ (.A1(_02266_),
    .A2(_03759_),
    .B1_N(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__mux2_2 _08855_ (.A0(\rvsingle.dp.rf.rf[20][24] ),
    .A1(\rvsingle.dp.rf.rf[21][24] ),
    .S(_01780_),
    .X(_03776_));
 sky130_fd_sc_hd__a21oi_2 _08856_ (.A1(_03776_),
    .A2(_01497_),
    .B1(_01565_),
    .Y(_03777_));
 sky130_fd_sc_hd__buf_1 _08857_ (.A(_01842_),
    .X(_03778_));
 sky130_fd_sc_hd__o21a_2 _08858_ (.A1(_01643_),
    .A2(\rvsingle.dp.rf.rf[22][24] ),
    .B1(_01648_),
    .X(_03779_));
 sky130_fd_sc_hd__o21ai_2 _08859_ (.A1(\rvsingle.dp.rf.rf[23][24] ),
    .A2(_03778_),
    .B1(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__mux4_2 _08860_ (.A0(\rvsingle.dp.rf.rf[16][24] ),
    .A1(\rvsingle.dp.rf.rf[17][24] ),
    .A2(\rvsingle.dp.rf.rf[18][24] ),
    .A3(\rvsingle.dp.rf.rf[19][24] ),
    .S0(_01493_),
    .S1(_01612_),
    .X(_03781_));
 sky130_fd_sc_hd__buf_1 _08861_ (.A(_01632_),
    .X(_03782_));
 sky130_fd_sc_hd__o2bb2ai_2 _08862_ (.A1_N(_03777_),
    .A2_N(_03780_),
    .B1(_03781_),
    .B2(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__mux4_2 _08863_ (.A0(\rvsingle.dp.rf.rf[24][24] ),
    .A1(\rvsingle.dp.rf.rf[25][24] ),
    .A2(\rvsingle.dp.rf.rf[26][24] ),
    .A3(\rvsingle.dp.rf.rf[27][24] ),
    .S0(_01137_),
    .S1(_01612_),
    .X(_03784_));
 sky130_fd_sc_hd__or2_2 _08864_ (.A(_01780_),
    .B(\rvsingle.dp.rf.rf[28][24] ),
    .X(_03785_));
 sky130_fd_sc_hd__o211a_2 _08865_ (.A1(\rvsingle.dp.rf.rf[29][24] ),
    .A2(_01540_),
    .B1(_01543_),
    .C1(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__mux2_2 _08866_ (.A0(\rvsingle.dp.rf.rf[30][24] ),
    .A1(\rvsingle.dp.rf.rf[31][24] ),
    .S(_01658_),
    .X(_03787_));
 sky130_fd_sc_hd__a21o_2 _08867_ (.A1(_01491_),
    .A2(_03787_),
    .B1(_01768_),
    .X(_03788_));
 sky130_fd_sc_hd__o221ai_2 _08868_ (.A1(_01512_),
    .A2(_03784_),
    .B1(_03786_),
    .B2(_03788_),
    .C1(_01506_),
    .Y(_03789_));
 sky130_fd_sc_hd__o211ai_2 _08869_ (.A1(_01117_),
    .A2(_03783_),
    .B1(_01682_),
    .C1(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__mux4_2 _08870_ (.A0(\rvsingle.dp.rf.rf[12][24] ),
    .A1(\rvsingle.dp.rf.rf[13][24] ),
    .A2(\rvsingle.dp.rf.rf[14][24] ),
    .A3(\rvsingle.dp.rf.rf[15][24] ),
    .S0(_01656_),
    .S1(_01260_),
    .X(_03791_));
 sky130_fd_sc_hd__nor2_2 _08871_ (.A(_02236_),
    .B(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__mux4_2 _08872_ (.A0(\rvsingle.dp.rf.rf[8][24] ),
    .A1(\rvsingle.dp.rf.rf[9][24] ),
    .A2(\rvsingle.dp.rf.rf[10][24] ),
    .A3(\rvsingle.dp.rf.rf[11][24] ),
    .S0(_01518_),
    .S1(_01626_),
    .X(_03793_));
 sky130_fd_sc_hd__o21ai_2 _08873_ (.A1(_03782_),
    .A2(_03793_),
    .B1(_01506_),
    .Y(_03794_));
 sky130_fd_sc_hd__mux4_2 _08874_ (.A0(\rvsingle.dp.rf.rf[4][24] ),
    .A1(\rvsingle.dp.rf.rf[5][24] ),
    .A2(\rvsingle.dp.rf.rf[6][24] ),
    .A3(\rvsingle.dp.rf.rf[7][24] ),
    .S0(_01562_),
    .S1(_01655_),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_2 _08875_ (.A0(\rvsingle.dp.rf.rf[0][24] ),
    .A1(\rvsingle.dp.rf.rf[1][24] ),
    .S(_02117_),
    .X(_03796_));
 sky130_fd_sc_hd__o21a_2 _08876_ (.A1(_01255_),
    .A2(\rvsingle.dp.rf.rf[2][24] ),
    .B1(_01530_),
    .X(_03797_));
 sky130_fd_sc_hd__o21a_2 _08877_ (.A1(_01677_),
    .A2(\rvsingle.dp.rf.rf[3][24] ),
    .B1(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__a211o_2 _08878_ (.A1(_03796_),
    .A2(_01543_),
    .B1(_01632_),
    .C1(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__o211ai_2 _08879_ (.A1(_02236_),
    .A2(_03795_),
    .B1(_03799_),
    .C1(_01157_),
    .Y(_03800_));
 sky130_fd_sc_hd__o211ai_2 _08880_ (.A1(_03792_),
    .A2(_03794_),
    .B1(_01378_),
    .C1(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__and4_2 _08881_ (.A(_01153_),
    .B(_03790_),
    .C(_03801_),
    .D(_01537_),
    .X(_03802_));
 sky130_fd_sc_hd__o21a_2 _08882_ (.A1(_01179_),
    .A2(_03802_),
    .B1(_01184_),
    .X(_03803_));
 sky130_fd_sc_hd__or2_2 _08883_ (.A(_01417_),
    .B(\rvsingle.dp.rf.rf[16][24] ),
    .X(_03804_));
 sky130_fd_sc_hd__o211ai_2 _08884_ (.A1(\rvsingle.dp.rf.rf[17][24] ),
    .A2(_01296_),
    .B1(_01717_),
    .C1(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__mux2_2 _08885_ (.A0(\rvsingle.dp.rf.rf[18][24] ),
    .A1(\rvsingle.dp.rf.rf[19][24] ),
    .S(_01192_),
    .X(_03806_));
 sky130_fd_sc_hd__a21oi_2 _08886_ (.A1(_01451_),
    .A2(_03806_),
    .B1(_01445_),
    .Y(_03807_));
 sky130_fd_sc_hd__mux4_2 _08887_ (.A0(\rvsingle.dp.rf.rf[20][24] ),
    .A1(\rvsingle.dp.rf.rf[21][24] ),
    .A2(\rvsingle.dp.rf.rf[22][24] ),
    .A3(\rvsingle.dp.rf.rf[23][24] ),
    .S0(_01469_),
    .S1(_01728_),
    .X(_03808_));
 sky130_fd_sc_hd__o2bb2a_2 _08888_ (.A1_N(_03805_),
    .A2_N(_03807_),
    .B1(_01722_),
    .B2(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__mux4_2 _08889_ (.A0(\rvsingle.dp.rf.rf[28][24] ),
    .A1(\rvsingle.dp.rf.rf[29][24] ),
    .A2(\rvsingle.dp.rf.rf[30][24] ),
    .A3(\rvsingle.dp.rf.rf[31][24] ),
    .S0(_01463_),
    .S1(_01471_),
    .X(_03810_));
 sky130_fd_sc_hd__mux4_2 _08890_ (.A0(\rvsingle.dp.rf.rf[24][24] ),
    .A1(\rvsingle.dp.rf.rf[25][24] ),
    .A2(\rvsingle.dp.rf.rf[26][24] ),
    .A3(\rvsingle.dp.rf.rf[27][24] ),
    .S0(_01328_),
    .S1(_01455_),
    .X(_03811_));
 sky130_fd_sc_hd__or2_2 _08891_ (.A(_01229_),
    .B(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__o211a_2 _08892_ (.A1(_01722_),
    .A2(_03810_),
    .B1(_01478_),
    .C1(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__a211o_2 _08893_ (.A1(_01219_),
    .A2(_03809_),
    .B1(_01316_),
    .C1(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__mux4_2 _08894_ (.A0(\rvsingle.dp.rf.rf[0][24] ),
    .A1(\rvsingle.dp.rf.rf[1][24] ),
    .A2(\rvsingle.dp.rf.rf[2][24] ),
    .A3(\rvsingle.dp.rf.rf[3][24] ),
    .S0(_01726_),
    .S1(_01728_),
    .X(_03815_));
 sky130_fd_sc_hd__mux4_2 _08895_ (.A0(\rvsingle.dp.rf.rf[4][24] ),
    .A1(\rvsingle.dp.rf.rf[5][24] ),
    .A2(\rvsingle.dp.rf.rf[6][24] ),
    .A3(\rvsingle.dp.rf.rf[7][24] ),
    .S0(_01726_),
    .S1(_01728_),
    .X(_03816_));
 sky130_fd_sc_hd__mux2_2 _08896_ (.A0(_03815_),
    .A1(_03816_),
    .S(_01445_),
    .X(_03817_));
 sky130_fd_sc_hd__mux4_2 _08897_ (.A0(\rvsingle.dp.rf.rf[8][24] ),
    .A1(\rvsingle.dp.rf.rf[9][24] ),
    .A2(\rvsingle.dp.rf.rf[10][24] ),
    .A3(\rvsingle.dp.rf.rf[11][24] ),
    .S0(_01463_),
    .S1(_01471_),
    .X(_03818_));
 sky130_fd_sc_hd__mux2_2 _08898_ (.A0(\rvsingle.dp.rf.rf[12][24] ),
    .A1(\rvsingle.dp.rf.rf[13][24] ),
    .S(_01335_),
    .X(_03819_));
 sky130_fd_sc_hd__or2_2 _08899_ (.A(_01828_),
    .B(\rvsingle.dp.rf.rf[14][24] ),
    .X(_03820_));
 sky130_fd_sc_hd__o211a_2 _08900_ (.A1(_02288_),
    .A2(\rvsingle.dp.rf.rf[15][24] ),
    .B1(_01433_),
    .C1(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__a211o_2 _08901_ (.A1(_03819_),
    .A2(_01437_),
    .B1(_01721_),
    .C1(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__o211a_2 _08902_ (.A1(_01703_),
    .A2(_03818_),
    .B1(_03822_),
    .C1(_01478_),
    .X(_03823_));
 sky130_fd_sc_hd__a211o_2 _08903_ (.A1(_01219_),
    .A2(_03817_),
    .B1(_03823_),
    .C1(_01450_),
    .X(_03824_));
 sky130_fd_sc_hd__and3_2 _08904_ (.A(_01248_),
    .B(_03814_),
    .C(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__or3_2 _08905_ (.A(_01184_),
    .B(_01179_),
    .C(_03802_),
    .X(_03826_));
 sky130_fd_sc_hd__nand3b_2 _08906_ (.A_N(_03803_),
    .B(_03825_),
    .C(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__a211oi_2 _08907_ (.A1(_01961_),
    .A2(Instr[31]),
    .B1(_01184_),
    .C1(_03802_),
    .Y(_03828_));
 sky130_fd_sc_hd__o21bai_2 _08908_ (.A1(_03828_),
    .A2(_03803_),
    .B1_N(_03825_),
    .Y(_03829_));
 sky130_fd_sc_hd__nand2_2 _08909_ (.A(_03827_),
    .B(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__inv_2 _08910_ (.A(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__o21a_2 _08911_ (.A1(_01848_),
    .A2(\rvsingle.dp.rf.rf[26][25] ),
    .B1(_01648_),
    .X(_03832_));
 sky130_fd_sc_hd__o21a_2 _08912_ (.A1(_03778_),
    .A2(\rvsingle.dp.rf.rf[27][25] ),
    .B1(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__or2b_2 _08913_ (.A(\rvsingle.dp.rf.rf[25][25] ),
    .B_N(_01126_),
    .X(_03834_));
 sky130_fd_sc_hd__o211a_2 _08914_ (.A1(_01257_),
    .A2(\rvsingle.dp.rf.rf[24][25] ),
    .B1(_03834_),
    .C1(_01856_),
    .X(_03835_));
 sky130_fd_sc_hd__nor2_2 _08915_ (.A(_01138_),
    .B(\rvsingle.dp.rf.rf[28][25] ),
    .Y(_03836_));
 sky130_fd_sc_hd__o21ai_2 _08916_ (.A1(\rvsingle.dp.rf.rf[29][25] ),
    .A2(_01488_),
    .B1(_01497_),
    .Y(_03837_));
 sky130_fd_sc_hd__nor2_2 _08917_ (.A(_01257_),
    .B(\rvsingle.dp.rf.rf[30][25] ),
    .Y(_03838_));
 sky130_fd_sc_hd__buf_1 _08918_ (.A(_01796_),
    .X(_03839_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08919_ (.A(_01531_),
    .X(_03840_));
 sky130_fd_sc_hd__o21ai_2 _08920_ (.A1(\rvsingle.dp.rf.rf[31][25] ),
    .A2(_03839_),
    .B1(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__o221ai_2 _08921_ (.A1(_03836_),
    .A2(_03837_),
    .B1(_03838_),
    .B2(_03841_),
    .C1(_03782_),
    .Y(_03842_));
 sky130_fd_sc_hd__o311ai_2 _08922_ (.A1(_03782_),
    .A2(_03833_),
    .A3(_03835_),
    .B1(_01117_),
    .C1(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__nor2_2 _08923_ (.A(_01138_),
    .B(\rvsingle.dp.rf.rf[20][25] ),
    .Y(_03844_));
 sky130_fd_sc_hd__and2b_2 _08924_ (.A_N(\rvsingle.dp.rf.rf[21][25] ),
    .B(_01643_),
    .X(_03845_));
 sky130_fd_sc_hd__nor2_2 _08925_ (.A(_01257_),
    .B(\rvsingle.dp.rf.rf[22][25] ),
    .Y(_03846_));
 sky130_fd_sc_hd__o21ai_2 _08926_ (.A1(\rvsingle.dp.rf.rf[23][25] ),
    .A2(_03839_),
    .B1(_03840_),
    .Y(_03847_));
 sky130_fd_sc_hd__o32ai_2 _08927_ (.A1(_01106_),
    .A2(_03844_),
    .A3(_03845_),
    .B1(_03846_),
    .B2(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__nor2_2 _08928_ (.A(_01257_),
    .B(\rvsingle.dp.rf.rf[18][25] ),
    .Y(_03849_));
 sky130_fd_sc_hd__o21ai_2 _08929_ (.A1(\rvsingle.dp.rf.rf[19][25] ),
    .A2(_03839_),
    .B1(_03840_),
    .Y(_03850_));
 sky130_fd_sc_hd__or2_2 _08930_ (.A(_01562_),
    .B(\rvsingle.dp.rf.rf[16][25] ),
    .X(_03851_));
 sky130_fd_sc_hd__o211ai_2 _08931_ (.A1(\rvsingle.dp.rf.rf[17][25] ),
    .A2(_03839_),
    .B1(_01497_),
    .C1(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__o211ai_2 _08932_ (.A1(_03849_),
    .A2(_03850_),
    .B1(_03852_),
    .C1(_02236_),
    .Y(_03853_));
 sky130_fd_sc_hd__o211ai_2 _08933_ (.A1(_01133_),
    .A2(_03848_),
    .B1(_03853_),
    .C1(_01157_),
    .Y(_03854_));
 sky130_fd_sc_hd__nand3_2 _08934_ (.A(_03843_),
    .B(_03854_),
    .C(_01147_),
    .Y(_03855_));
 sky130_fd_sc_hd__nor2_2 _08935_ (.A(_01127_),
    .B(\rvsingle.dp.rf.rf[2][25] ),
    .Y(_03856_));
 sky130_fd_sc_hd__buf_1 _08936_ (.A(_01646_),
    .X(_03857_));
 sky130_fd_sc_hd__o21ai_2 _08937_ (.A1(\rvsingle.dp.rf.rf[3][25] ),
    .A2(_03857_),
    .B1(_03840_),
    .Y(_03858_));
 sky130_fd_sc_hd__nor2_2 _08938_ (.A(_01127_),
    .B(\rvsingle.dp.rf.rf[0][25] ),
    .Y(_03859_));
 sky130_fd_sc_hd__o21ai_2 _08939_ (.A1(\rvsingle.dp.rf.rf[1][25] ),
    .A2(_03778_),
    .B1(_01856_),
    .Y(_03860_));
 sky130_fd_sc_hd__o221a_2 _08940_ (.A1(_03856_),
    .A2(_03858_),
    .B1(_03859_),
    .B2(_03860_),
    .C1(_02236_),
    .X(_03861_));
 sky130_fd_sc_hd__or2_2 _08941_ (.A(_01643_),
    .B(\rvsingle.dp.rf.rf[6][25] ),
    .X(_03862_));
 sky130_fd_sc_hd__o211ai_2 _08942_ (.A1(_03778_),
    .A2(\rvsingle.dp.rf.rf[7][25] ),
    .B1(_01106_),
    .C1(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__o21ba_2 _08943_ (.A1(_01098_),
    .A2(\rvsingle.dp.rf.rf[4][25] ),
    .B1_N(_01105_),
    .X(_03864_));
 sky130_fd_sc_hd__o21ai_2 _08944_ (.A1(_03778_),
    .A2(\rvsingle.dp.rf.rf[5][25] ),
    .B1(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__a31o_2 _08945_ (.A1(_03863_),
    .A2(_03782_),
    .A3(_03865_),
    .B1(_01506_),
    .X(_03866_));
 sky130_fd_sc_hd__nor2_2 _08946_ (.A(_01127_),
    .B(\rvsingle.dp.rf.rf[10][25] ),
    .Y(_03867_));
 sky130_fd_sc_hd__o21ai_2 _08947_ (.A1(\rvsingle.dp.rf.rf[11][25] ),
    .A2(_03857_),
    .B1(_03840_),
    .Y(_03868_));
 sky130_fd_sc_hd__or2b_2 _08948_ (.A(\rvsingle.dp.rf.rf[9][25] ),
    .B_N(_01126_),
    .X(_03869_));
 sky130_fd_sc_hd__o211ai_2 _08949_ (.A1(_01257_),
    .A2(\rvsingle.dp.rf.rf[8][25] ),
    .B1(_03869_),
    .C1(_01856_),
    .Y(_03870_));
 sky130_fd_sc_hd__o21ai_2 _08950_ (.A1(_03867_),
    .A2(_03868_),
    .B1(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__nor2_2 _08951_ (.A(_01257_),
    .B(\rvsingle.dp.rf.rf[12][25] ),
    .Y(_03872_));
 sky130_fd_sc_hd__o21ai_2 _08952_ (.A1(\rvsingle.dp.rf.rf[13][25] ),
    .A2(_03857_),
    .B1(_01856_),
    .Y(_03873_));
 sky130_fd_sc_hd__o21a_2 _08953_ (.A1(_01666_),
    .A2(\rvsingle.dp.rf.rf[14][25] ),
    .B1(_01612_),
    .X(_03874_));
 sky130_fd_sc_hd__o21ai_2 _08954_ (.A1(\rvsingle.dp.rf.rf[15][25] ),
    .A2(_03778_),
    .B1(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__o211ai_2 _08955_ (.A1(_03872_),
    .A2(_03873_),
    .B1(_03782_),
    .C1(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__o211ai_2 _08956_ (.A1(_01113_),
    .A2(_03871_),
    .B1(_03876_),
    .C1(_01117_),
    .Y(_03877_));
 sky130_fd_sc_hd__o211ai_2 _08957_ (.A1(_03861_),
    .A2(_03866_),
    .B1(_01378_),
    .C1(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__o211a_2 _08958_ (.A1(_02212_),
    .A2(_01962_),
    .B1(_03855_),
    .C1(_03878_),
    .X(WriteData[25]));
 sky130_fd_sc_hd__nand2_2 _08959_ (.A(_01085_),
    .B(WriteData[25]),
    .Y(_03879_));
 sky130_fd_sc_hd__a21oi_2 _08960_ (.A1(_01581_),
    .A2(_03879_),
    .B1(_01837_),
    .Y(_03880_));
 sky130_fd_sc_hd__and3_2 _08961_ (.A(_01837_),
    .B(_01581_),
    .C(_03879_),
    .X(_03881_));
 sky130_fd_sc_hd__mux4_2 _08962_ (.A0(\rvsingle.dp.rf.rf[20][25] ),
    .A1(\rvsingle.dp.rf.rf[21][25] ),
    .A2(\rvsingle.dp.rf.rf[22][25] ),
    .A3(\rvsingle.dp.rf.rf[23][25] ),
    .S0(_01194_),
    .S1(_01201_),
    .X(_03882_));
 sky130_fd_sc_hd__nor2_2 _08963_ (.A(_01209_),
    .B(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__mux2_2 _08964_ (.A0(\rvsingle.dp.rf.rf[16][25] ),
    .A1(\rvsingle.dp.rf.rf[17][25] ),
    .S(_01194_),
    .X(_03884_));
 sky130_fd_sc_hd__or2_2 _08965_ (.A(_01194_),
    .B(\rvsingle.dp.rf.rf[18][25] ),
    .X(_03885_));
 sky130_fd_sc_hd__o211a_2 _08966_ (.A1(_01298_),
    .A2(\rvsingle.dp.rf.rf[19][25] ),
    .B1(_01303_),
    .C1(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__a211oi_2 _08967_ (.A1(_03884_),
    .A2(_01311_),
    .B1(_01231_),
    .C1(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__mux4_2 _08968_ (.A0(\rvsingle.dp.rf.rf[28][25] ),
    .A1(\rvsingle.dp.rf.rf[29][25] ),
    .A2(\rvsingle.dp.rf.rf[30][25] ),
    .A3(\rvsingle.dp.rf.rf[31][25] ),
    .S0(_01194_),
    .S1(_01303_),
    .X(_03888_));
 sky130_fd_sc_hd__mux4_2 _08969_ (.A0(\rvsingle.dp.rf.rf[24][25] ),
    .A1(\rvsingle.dp.rf.rf[25][25] ),
    .A2(\rvsingle.dp.rf.rf[26][25] ),
    .A3(\rvsingle.dp.rf.rf[27][25] ),
    .S0(_01330_),
    .S1(_01302_),
    .X(_03889_));
 sky130_fd_sc_hd__o21a_2 _08970_ (.A1(_01231_),
    .A2(_03889_),
    .B1(_01223_),
    .X(_03890_));
 sky130_fd_sc_hd__o21ai_2 _08971_ (.A1(_01209_),
    .A2(_03888_),
    .B1(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__o311ai_2 _08972_ (.A1(_01223_),
    .A2(_03883_),
    .A3(_03887_),
    .B1(_01189_),
    .C1(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__mux4_2 _08973_ (.A0(\rvsingle.dp.rf.rf[8][25] ),
    .A1(\rvsingle.dp.rf.rf[9][25] ),
    .A2(\rvsingle.dp.rf.rf[10][25] ),
    .A3(\rvsingle.dp.rf.rf[11][25] ),
    .S0(_01330_),
    .S1(_01302_),
    .X(_03893_));
 sky130_fd_sc_hd__or2_2 _08974_ (.A(_01193_),
    .B(\rvsingle.dp.rf.rf[12][25] ),
    .X(_03894_));
 sky130_fd_sc_hd__o211ai_2 _08975_ (.A1(\rvsingle.dp.rf.rf[13][25] ),
    .A2(_01297_),
    .B1(_01310_),
    .C1(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__o21a_2 _08976_ (.A1(_01193_),
    .A2(\rvsingle.dp.rf.rf[14][25] ),
    .B1(_01200_),
    .X(_03896_));
 sky130_fd_sc_hd__o21ai_2 _08977_ (.A1(\rvsingle.dp.rf.rf[15][25] ),
    .A2(_01297_),
    .B1(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand3_2 _08978_ (.A(_03895_),
    .B(_01915_),
    .C(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__o211a_2 _08979_ (.A1(_01915_),
    .A2(_03893_),
    .B1(_03898_),
    .C1(_01222_),
    .X(_03899_));
 sky130_fd_sc_hd__mux4_2 _08980_ (.A0(\rvsingle.dp.rf.rf[4][25] ),
    .A1(\rvsingle.dp.rf.rf[5][25] ),
    .A2(\rvsingle.dp.rf.rf[6][25] ),
    .A3(\rvsingle.dp.rf.rf[7][25] ),
    .S0(_01330_),
    .S1(_01302_),
    .X(_03900_));
 sky130_fd_sc_hd__mux2_2 _08981_ (.A0(\rvsingle.dp.rf.rf[0][25] ),
    .A1(\rvsingle.dp.rf.rf[1][25] ),
    .S(_01336_),
    .X(_03901_));
 sky130_fd_sc_hd__or2_2 _08982_ (.A(_01463_),
    .B(\rvsingle.dp.rf.rf[2][25] ),
    .X(_03902_));
 sky130_fd_sc_hd__o211a_2 _08983_ (.A1(_01296_),
    .A2(\rvsingle.dp.rf.rf[3][25] ),
    .B1(_01434_),
    .C1(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__a211o_2 _08984_ (.A1(_03901_),
    .A2(_01310_),
    .B1(_01230_),
    .C1(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__o211a_2 _08985_ (.A1(_02191_),
    .A2(_03900_),
    .B1(_03904_),
    .C1(_01219_),
    .X(_03905_));
 sky130_fd_sc_hd__or3_2 _08986_ (.A(_01189_),
    .B(_03899_),
    .C(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__o211ai_2 _08987_ (.A1(_01351_),
    .A2(_01203_),
    .B1(_03892_),
    .C1(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__o21ai_2 _08988_ (.A1(_03880_),
    .A2(_03881_),
    .B1(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__or3_2 _08989_ (.A(_03907_),
    .B(_03880_),
    .C(_03881_),
    .X(_03909_));
 sky130_fd_sc_hd__and3_2 _08990_ (.A(_03831_),
    .B(_03908_),
    .C(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__mux4_2 _08991_ (.A0(\rvsingle.dp.rf.rf[24][27] ),
    .A1(\rvsingle.dp.rf.rf[25][27] ),
    .A2(\rvsingle.dp.rf.rf[26][27] ),
    .A3(\rvsingle.dp.rf.rf[27][27] ),
    .S0(_01330_),
    .S1(_01302_),
    .X(_03911_));
 sky130_fd_sc_hd__mux2_2 _08992_ (.A0(\rvsingle.dp.rf.rf[28][27] ),
    .A1(\rvsingle.dp.rf.rf[29][27] ),
    .S(_01193_),
    .X(_03912_));
 sky130_fd_sc_hd__or2_2 _08993_ (.A(_01432_),
    .B(\rvsingle.dp.rf.rf[30][27] ),
    .X(_03913_));
 sky130_fd_sc_hd__o211a_2 _08994_ (.A1(_01296_),
    .A2(\rvsingle.dp.rf.rf[31][27] ),
    .B1(_01200_),
    .C1(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__a211o_2 _08995_ (.A1(_03912_),
    .A2(_01310_),
    .B1(_02191_),
    .C1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__o211ai_2 _08996_ (.A1(_01231_),
    .A2(_03911_),
    .B1(_03915_),
    .C1(_01223_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand2_2 _08997_ (.A(_03916_),
    .B(_01189_),
    .Y(_03917_));
 sky130_fd_sc_hd__mux4_2 _08998_ (.A0(\rvsingle.dp.rf.rf[20][27] ),
    .A1(\rvsingle.dp.rf.rf[21][27] ),
    .A2(\rvsingle.dp.rf.rf[22][27] ),
    .A3(\rvsingle.dp.rf.rf[23][27] ),
    .S0(_01337_),
    .S1(_01201_),
    .X(_03918_));
 sky130_fd_sc_hd__mux2_2 _08999_ (.A0(\rvsingle.dp.rf.rf[16][27] ),
    .A1(\rvsingle.dp.rf.rf[17][27] ),
    .S(_01193_),
    .X(_03919_));
 sky130_fd_sc_hd__or2_2 _09000_ (.A(_01242_),
    .B(\rvsingle.dp.rf.rf[18][27] ),
    .X(_03920_));
 sky130_fd_sc_hd__o211a_2 _09001_ (.A1(_01943_),
    .A2(\rvsingle.dp.rf.rf[19][27] ),
    .B1(_01451_),
    .C1(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__a211o_2 _09002_ (.A1(_03919_),
    .A2(_01310_),
    .B1(_01915_),
    .C1(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__o211a_2 _09003_ (.A1(_01209_),
    .A2(_03918_),
    .B1(_03922_),
    .C1(_01219_),
    .X(_03923_));
 sky130_fd_sc_hd__inv_2 _09004_ (.A(net212),
    .Y(_03924_));
 sky130_fd_sc_hd__nor2_2 _09005_ (.A(_01193_),
    .B(\rvsingle.dp.rf.rf[8][27] ),
    .Y(_03925_));
 sky130_fd_sc_hd__a211o_2 _09006_ (.A1(_03924_),
    .A2(_01330_),
    .B1(_01451_),
    .C1(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__mux2_2 _09007_ (.A0(\rvsingle.dp.rf.rf[10][27] ),
    .A1(\rvsingle.dp.rf.rf[11][27] ),
    .S(_01242_),
    .X(_03927_));
 sky130_fd_sc_hd__a21oi_2 _09008_ (.A1(_01302_),
    .A2(_03927_),
    .B1(_01230_),
    .Y(_03928_));
 sky130_fd_sc_hd__mux4_2 _09009_ (.A0(\rvsingle.dp.rf.rf[12][27] ),
    .A1(\rvsingle.dp.rf.rf[13][27] ),
    .A2(\rvsingle.dp.rf.rf[14][27] ),
    .A3(\rvsingle.dp.rf.rf[15][27] ),
    .S0(_01336_),
    .S1(_01200_),
    .X(_03929_));
 sky130_fd_sc_hd__o2bb2a_2 _09010_ (.A1_N(_03926_),
    .A2_N(_03928_),
    .B1(_02191_),
    .B2(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__mux4_2 _09011_ (.A0(\rvsingle.dp.rf.rf[4][27] ),
    .A1(\rvsingle.dp.rf.rf[5][27] ),
    .A2(\rvsingle.dp.rf.rf[6][27] ),
    .A3(\rvsingle.dp.rf.rf[7][27] ),
    .S0(_01336_),
    .S1(_01451_),
    .X(_03931_));
 sky130_fd_sc_hd__or2_2 _09012_ (.A(_01192_),
    .B(\rvsingle.dp.rf.rf[0][27] ),
    .X(_03932_));
 sky130_fd_sc_hd__o211ai_2 _09013_ (.A1(\rvsingle.dp.rf.rf[1][27] ),
    .A2(_01441_),
    .B1(_01437_),
    .C1(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__or2_2 _09014_ (.A(_01192_),
    .B(\rvsingle.dp.rf.rf[2][27] ),
    .X(_03934_));
 sky130_fd_sc_hd__o211ai_2 _09015_ (.A1(_01441_),
    .A2(\rvsingle.dp.rf.rf[3][27] ),
    .B1(_01434_),
    .C1(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__a31o_2 _09016_ (.A1(_01461_),
    .A2(_03933_),
    .A3(_03935_),
    .B1(_01447_),
    .X(_03936_));
 sky130_fd_sc_hd__o21ba_2 _09017_ (.A1(_02191_),
    .A2(_03931_),
    .B1_N(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__a211o_2 _09018_ (.A1(_03930_),
    .A2(_01223_),
    .B1(_01189_),
    .C1(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__o211ai_2 _09019_ (.A1(_03917_),
    .A2(_03923_),
    .B1(_01248_),
    .C1(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__mux2_2 _09020_ (.A0(\rvsingle.dp.rf.rf[16][27] ),
    .A1(\rvsingle.dp.rf.rf[17][27] ),
    .S(_01269_),
    .X(_03940_));
 sky130_fd_sc_hd__o21a_2 _09021_ (.A1(_01098_),
    .A2(\rvsingle.dp.rf.rf[18][27] ),
    .B1(_01626_),
    .X(_03941_));
 sky130_fd_sc_hd__o21a_2 _09022_ (.A1(_01089_),
    .A2(\rvsingle.dp.rf.rf[19][27] ),
    .B1(_03941_),
    .X(_03942_));
 sky130_fd_sc_hd__a211oi_2 _09023_ (.A1(_03940_),
    .A2(_01093_),
    .B1(_01113_),
    .C1(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__or2_2 _09024_ (.A(_01643_),
    .B(\rvsingle.dp.rf.rf[20][27] ),
    .X(_03944_));
 sky130_fd_sc_hd__o211ai_2 _09025_ (.A1(\rvsingle.dp.rf.rf[21][27] ),
    .A2(_01089_),
    .B1(_01093_),
    .C1(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__o21a_2 _09026_ (.A1(_01098_),
    .A2(\rvsingle.dp.rf.rf[22][27] ),
    .B1(_01655_),
    .X(_03946_));
 sky130_fd_sc_hd__o21ai_2 _09027_ (.A1(\rvsingle.dp.rf.rf[23][27] ),
    .A2(_01089_),
    .B1(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__a31o_2 _09028_ (.A1(_03945_),
    .A2(_03782_),
    .A3(_03947_),
    .B1(_01506_),
    .X(_03948_));
 sky130_fd_sc_hd__mux4_2 _09029_ (.A0(\rvsingle.dp.rf.rf[28][27] ),
    .A1(\rvsingle.dp.rf.rf[29][27] ),
    .A2(\rvsingle.dp.rf.rf[30][27] ),
    .A3(\rvsingle.dp.rf.rf[31][27] ),
    .S0(_01559_),
    .S1(_03840_),
    .X(_03949_));
 sky130_fd_sc_hd__or2_2 _09030_ (.A(_01256_),
    .B(\rvsingle.dp.rf.rf[24][27] ),
    .X(_03950_));
 sky130_fd_sc_hd__o21ai_2 _09031_ (.A1(_03839_),
    .A2(\rvsingle.dp.rf.rf[25][27] ),
    .B1(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__or2_2 _09032_ (.A(_01256_),
    .B(\rvsingle.dp.rf.rf[26][27] ),
    .X(_03952_));
 sky130_fd_sc_hd__o211ai_2 _09033_ (.A1(_03839_),
    .A2(\rvsingle.dp.rf.rf[27][27] ),
    .B1(_03840_),
    .C1(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__o211ai_2 _09034_ (.A1(_01106_),
    .A2(_03951_),
    .B1(_03953_),
    .C1(_02236_),
    .Y(_03954_));
 sky130_fd_sc_hd__o211ai_2 _09035_ (.A1(_01133_),
    .A2(_03949_),
    .B1(_03954_),
    .C1(_01117_),
    .Y(_03955_));
 sky130_fd_sc_hd__o211ai_2 _09036_ (.A1(_03943_),
    .A2(_03948_),
    .B1(_01147_),
    .C1(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__o21ba_2 _09037_ (.A1(_01848_),
    .A2(\rvsingle.dp.rf.rf[0][27] ),
    .B1_N(_01605_),
    .X(_03957_));
 sky130_fd_sc_hd__o21ai_2 _09038_ (.A1(_03857_),
    .A2(\rvsingle.dp.rf.rf[1][27] ),
    .B1(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__o21a_2 _09039_ (.A1(_01848_),
    .A2(\rvsingle.dp.rf.rf[2][27] ),
    .B1(_01612_),
    .X(_03959_));
 sky130_fd_sc_hd__o21ai_2 _09040_ (.A1(\rvsingle.dp.rf.rf[3][27] ),
    .A2(_03778_),
    .B1(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__and3_2 _09041_ (.A(_02236_),
    .B(_03958_),
    .C(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__or2_2 _09042_ (.A(_01643_),
    .B(\rvsingle.dp.rf.rf[4][27] ),
    .X(_03962_));
 sky130_fd_sc_hd__o211ai_2 _09043_ (.A1(\rvsingle.dp.rf.rf[5][27] ),
    .A2(_03778_),
    .B1(_01093_),
    .C1(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__or2_2 _09044_ (.A(_01744_),
    .B(\rvsingle.dp.rf.rf[6][27] ),
    .X(_03964_));
 sky130_fd_sc_hd__o211ai_2 _09045_ (.A1(_03857_),
    .A2(\rvsingle.dp.rf.rf[7][27] ),
    .B1(_01106_),
    .C1(_03964_),
    .Y(_03965_));
 sky130_fd_sc_hd__a31o_2 _09046_ (.A1(_03963_),
    .A2(_03965_),
    .A3(_03782_),
    .B1(_01506_),
    .X(_03966_));
 sky130_fd_sc_hd__o21a_2 _09047_ (.A1(_01744_),
    .A2(\rvsingle.dp.rf.rf[10][27] ),
    .B1(_01105_),
    .X(_03967_));
 sky130_fd_sc_hd__o21a_2 _09048_ (.A1(_03857_),
    .A2(\rvsingle.dp.rf.rf[11][27] ),
    .B1(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__nor2_2 _09049_ (.A(_01138_),
    .B(\rvsingle.dp.rf.rf[8][27] ),
    .Y(_03969_));
 sky130_fd_sc_hd__a211oi_2 _09050_ (.A1(_03924_),
    .A2(_01127_),
    .B1(_01106_),
    .C1(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__or2_2 _09051_ (.A(_01603_),
    .B(\rvsingle.dp.rf.rf[12][27] ),
    .X(_03971_));
 sky130_fd_sc_hd__o211ai_2 _09052_ (.A1(\rvsingle.dp.rf.rf[13][27] ),
    .A2(_03857_),
    .B1(_01856_),
    .C1(_03971_),
    .Y(_03972_));
 sky130_fd_sc_hd__o21a_2 _09053_ (.A1(_01744_),
    .A2(\rvsingle.dp.rf.rf[14][27] ),
    .B1(_01648_),
    .X(_03973_));
 sky130_fd_sc_hd__o21ai_2 _09054_ (.A1(\rvsingle.dp.rf.rf[15][27] ),
    .A2(_03857_),
    .B1(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand3_2 _09055_ (.A(_03972_),
    .B(_01512_),
    .C(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__o311ai_2 _09056_ (.A1(_03782_),
    .A2(_03968_),
    .A3(_03970_),
    .B1(_01117_),
    .C1(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__o211ai_2 _09057_ (.A1(_03961_),
    .A2(_03966_),
    .B1(_03976_),
    .C1(_01378_),
    .Y(_03977_));
 sky130_fd_sc_hd__a41o_2 _09058_ (.A1(_01153_),
    .A2(_03956_),
    .A3(_03977_),
    .A4(_01482_),
    .B1(_01184_),
    .X(_03978_));
 sky130_fd_sc_hd__a21oi_2 _09059_ (.A1(Instr[31]),
    .A2(_01961_),
    .B1(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__and4_2 _09060_ (.A(_01153_),
    .B(_03956_),
    .C(_03977_),
    .D(_01084_),
    .X(_03980_));
 sky130_fd_sc_hd__o21a_2 _09061_ (.A1(_01180_),
    .A2(_03980_),
    .B1(_01184_),
    .X(_03981_));
 sky130_fd_sc_hd__nor3_2 _09062_ (.A(_03939_),
    .B(_03979_),
    .C(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__o21ai_2 _09063_ (.A1(_03979_),
    .A2(_03981_),
    .B1(_03939_),
    .Y(_03983_));
 sky130_fd_sc_hd__or2b_2 _09064_ (.A(_03982_),
    .B_N(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__o21a_2 _09065_ (.A1(\rvsingle.dp.rf.rf[3][26] ),
    .A2(_01297_),
    .B1(_01302_),
    .X(_03985_));
 sky130_fd_sc_hd__or2_2 _09066_ (.A(_01337_),
    .B(\rvsingle.dp.rf.rf[2][26] ),
    .X(_03986_));
 sky130_fd_sc_hd__mux2_2 _09067_ (.A0(\rvsingle.dp.rf.rf[0][26] ),
    .A1(\rvsingle.dp.rf.rf[1][26] ),
    .S(_01337_),
    .X(_03987_));
 sky130_fd_sc_hd__a221oi_2 _09068_ (.A1(_03985_),
    .A2(_03986_),
    .B1(_03987_),
    .B2(_01310_),
    .C1(_01915_),
    .Y(_03988_));
 sky130_fd_sc_hd__mux2_2 _09069_ (.A0(\rvsingle.dp.rf.rf[4][26] ),
    .A1(\rvsingle.dp.rf.rf[5][26] ),
    .S(_01337_),
    .X(_03989_));
 sky130_fd_sc_hd__or2_2 _09070_ (.A(_01330_),
    .B(\rvsingle.dp.rf.rf[6][26] ),
    .X(_03990_));
 sky130_fd_sc_hd__o211a_2 _09071_ (.A1(_01297_),
    .A2(\rvsingle.dp.rf.rf[7][26] ),
    .B1(_01201_),
    .C1(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__a211oi_2 _09072_ (.A1(_03989_),
    .A2(_01310_),
    .B1(_01209_),
    .C1(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__o21a_2 _09073_ (.A1(\rvsingle.dp.rf.rf[11][26] ),
    .A2(_01943_),
    .B1(_01451_),
    .X(_03993_));
 sky130_fd_sc_hd__o21ai_2 _09074_ (.A1(_01194_),
    .A2(\rvsingle.dp.rf.rf[10][26] ),
    .B1(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__or2_2 _09075_ (.A(_01330_),
    .B(\rvsingle.dp.rf.rf[8][26] ),
    .X(_03995_));
 sky130_fd_sc_hd__o211ai_2 _09076_ (.A1(\rvsingle.dp.rf.rf[9][26] ),
    .A2(_01297_),
    .B1(_01310_),
    .C1(_03995_),
    .Y(_03996_));
 sky130_fd_sc_hd__mux2_2 _09077_ (.A0(\rvsingle.dp.rf.rf[12][26] ),
    .A1(\rvsingle.dp.rf.rf[13][26] ),
    .S(_01193_),
    .X(_03997_));
 sky130_fd_sc_hd__or2_2 _09078_ (.A(_01432_),
    .B(\rvsingle.dp.rf.rf[14][26] ),
    .X(_03998_));
 sky130_fd_sc_hd__o211a_2 _09079_ (.A1(_01943_),
    .A2(\rvsingle.dp.rf.rf[15][26] ),
    .B1(_01200_),
    .C1(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__a211oi_2 _09080_ (.A1(_03997_),
    .A2(_01310_),
    .B1(_02191_),
    .C1(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__a311o_2 _09081_ (.A1(_02191_),
    .A2(_03994_),
    .A3(_03996_),
    .B1(_01219_),
    .C1(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__o311a_2 _09082_ (.A1(_01223_),
    .A2(_03988_),
    .A3(_03992_),
    .B1(_01317_),
    .C1(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__mux4_2 _09083_ (.A0(\rvsingle.dp.rf.rf[28][26] ),
    .A1(\rvsingle.dp.rf.rf[29][26] ),
    .A2(\rvsingle.dp.rf.rf[30][26] ),
    .A3(\rvsingle.dp.rf.rf[31][26] ),
    .S0(_01330_),
    .S1(_01302_),
    .X(_04003_));
 sky130_fd_sc_hd__mux2_2 _09084_ (.A0(\rvsingle.dp.rf.rf[26][26] ),
    .A1(\rvsingle.dp.rf.rf[27][26] ),
    .S(_01193_),
    .X(_04004_));
 sky130_fd_sc_hd__or2_2 _09085_ (.A(_01432_),
    .B(\rvsingle.dp.rf.rf[24][26] ),
    .X(_04005_));
 sky130_fd_sc_hd__o211a_2 _09086_ (.A1(\rvsingle.dp.rf.rf[25][26] ),
    .A2(_01943_),
    .B1(_01717_),
    .C1(_04005_),
    .X(_04006_));
 sky130_fd_sc_hd__a211o_2 _09087_ (.A1(_01201_),
    .A2(_04004_),
    .B1(_04006_),
    .C1(_01915_),
    .X(_04007_));
 sky130_fd_sc_hd__o211ai_2 _09088_ (.A1(_01209_),
    .A2(_04003_),
    .B1(_01223_),
    .C1(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__mux4_2 _09089_ (.A0(\rvsingle.dp.rf.rf[16][26] ),
    .A1(\rvsingle.dp.rf.rf[17][26] ),
    .A2(\rvsingle.dp.rf.rf[18][26] ),
    .A3(\rvsingle.dp.rf.rf[19][26] ),
    .S0(_01337_),
    .S1(_01302_),
    .X(_04009_));
 sky130_fd_sc_hd__mux4_2 _09090_ (.A0(\rvsingle.dp.rf.rf[20][26] ),
    .A1(\rvsingle.dp.rf.rf[21][26] ),
    .A2(\rvsingle.dp.rf.rf[22][26] ),
    .A3(\rvsingle.dp.rf.rf[23][26] ),
    .S0(_01242_),
    .S1(_01200_),
    .X(_04010_));
 sky130_fd_sc_hd__o21ai_2 _09091_ (.A1(_02191_),
    .A2(_04010_),
    .B1(_01218_),
    .Y(_04011_));
 sky130_fd_sc_hd__o21bai_2 _09092_ (.A1(_01231_),
    .A2(_04009_),
    .B1_N(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__a31o_2 _09093_ (.A1(_04008_),
    .A2(_04012_),
    .A3(_01189_),
    .B1(_02469_),
    .X(_04013_));
 sky130_fd_sc_hd__mux2_2 _09094_ (.A0(\rvsingle.dp.rf.rf[0][26] ),
    .A1(\rvsingle.dp.rf.rf[1][26] ),
    .S(_01269_),
    .X(_04014_));
 sky130_fd_sc_hd__or2_2 _09095_ (.A(_01126_),
    .B(\rvsingle.dp.rf.rf[2][26] ),
    .X(_04015_));
 sky130_fd_sc_hd__o211a_2 _09096_ (.A1(_03857_),
    .A2(\rvsingle.dp.rf.rf[3][26] ),
    .B1(_03840_),
    .C1(_04015_),
    .X(_04016_));
 sky130_fd_sc_hd__a211oi_2 _09097_ (.A1(_04014_),
    .A2(_01093_),
    .B1(_03782_),
    .C1(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__inv_2 _09098_ (.A(\rvsingle.dp.rf.rf[7][26] ),
    .Y(_04018_));
 sky130_fd_sc_hd__o21ai_2 _09099_ (.A1(_01138_),
    .A2(\rvsingle.dp.rf.rf[6][26] ),
    .B1(_03840_),
    .Y(_04019_));
 sky130_fd_sc_hd__a21oi_2 _09100_ (.A1(_04018_),
    .A2(_01099_),
    .B1(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__or2_2 _09101_ (.A(_01603_),
    .B(\rvsingle.dp.rf.rf[4][26] ),
    .X(_04021_));
 sky130_fd_sc_hd__o211a_2 _09102_ (.A1(\rvsingle.dp.rf.rf[5][26] ),
    .A2(_03839_),
    .B1(_01856_),
    .C1(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__o31ai_2 _09103_ (.A1(_02236_),
    .A2(_04020_),
    .A3(_04022_),
    .B1(_01157_),
    .Y(_04023_));
 sky130_fd_sc_hd__mux4_2 _09104_ (.A0(\rvsingle.dp.rf.rf[12][26] ),
    .A1(\rvsingle.dp.rf.rf[13][26] ),
    .A2(\rvsingle.dp.rf.rf[14][26] ),
    .A3(\rvsingle.dp.rf.rf[15][26] ),
    .S0(_01098_),
    .S1(_03840_),
    .X(_04024_));
 sky130_fd_sc_hd__nor2_2 _09105_ (.A(_01257_),
    .B(\rvsingle.dp.rf.rf[8][26] ),
    .Y(_04025_));
 sky130_fd_sc_hd__o21ai_2 _09106_ (.A1(\rvsingle.dp.rf.rf[9][26] ),
    .A2(_03857_),
    .B1(_01856_),
    .Y(_04026_));
 sky130_fd_sc_hd__o21a_2 _09107_ (.A1(_01848_),
    .A2(\rvsingle.dp.rf.rf[10][26] ),
    .B1(_01612_),
    .X(_04027_));
 sky130_fd_sc_hd__o21ai_2 _09108_ (.A1(\rvsingle.dp.rf.rf[11][26] ),
    .A2(_03778_),
    .B1(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__o211ai_2 _09109_ (.A1(_04025_),
    .A2(_04026_),
    .B1(_02236_),
    .C1(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__o211ai_2 _09110_ (.A1(_01133_),
    .A2(_04024_),
    .B1(_04029_),
    .C1(_01117_),
    .Y(_04030_));
 sky130_fd_sc_hd__o211ai_2 _09111_ (.A1(_04017_),
    .A2(_04023_),
    .B1(_01378_),
    .C1(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__o21ba_2 _09112_ (.A1(_01126_),
    .A2(\rvsingle.dp.rf.rf[20][26] ),
    .B1_N(_01531_),
    .X(_04032_));
 sky130_fd_sc_hd__o21ai_2 _09113_ (.A1(_03839_),
    .A2(\rvsingle.dp.rf.rf[21][26] ),
    .B1(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__o21a_2 _09114_ (.A1(_01126_),
    .A2(\rvsingle.dp.rf.rf[22][26] ),
    .B1(_01605_),
    .X(_04034_));
 sky130_fd_sc_hd__o21ai_2 _09115_ (.A1(\rvsingle.dp.rf.rf[23][26] ),
    .A2(_03839_),
    .B1(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__and3_2 _09116_ (.A(_04033_),
    .B(_04035_),
    .C(_01512_),
    .X(_04036_));
 sky130_fd_sc_hd__nor2_2 _09117_ (.A(_01127_),
    .B(\rvsingle.dp.rf.rf[16][26] ),
    .Y(_04037_));
 sky130_fd_sc_hd__o21ai_2 _09118_ (.A1(\rvsingle.dp.rf.rf[17][26] ),
    .A2(_03839_),
    .B1(_01856_),
    .Y(_04038_));
 sky130_fd_sc_hd__o21a_2 _09119_ (.A1(_01666_),
    .A2(\rvsingle.dp.rf.rf[18][26] ),
    .B1(_01626_),
    .X(_04039_));
 sky130_fd_sc_hd__o21ai_2 _09120_ (.A1(\rvsingle.dp.rf.rf[19][26] ),
    .A2(_03778_),
    .B1(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__o211a_2 _09121_ (.A1(_04037_),
    .A2(_04038_),
    .B1(_01132_),
    .C1(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__mux4_2 _09122_ (.A0(\rvsingle.dp.rf.rf[28][26] ),
    .A1(\rvsingle.dp.rf.rf[29][26] ),
    .A2(\rvsingle.dp.rf.rf[30][26] ),
    .A3(\rvsingle.dp.rf.rf[31][26] ),
    .S0(_01643_),
    .S1(_01491_),
    .X(_04042_));
 sky130_fd_sc_hd__or2_2 _09123_ (.A(_01614_),
    .B(\rvsingle.dp.rf.rf[24][26] ),
    .X(_04043_));
 sky130_fd_sc_hd__o21ai_2 _09124_ (.A1(_01488_),
    .A2(\rvsingle.dp.rf.rf[25][26] ),
    .B1(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__or2_2 _09125_ (.A(_01614_),
    .B(\rvsingle.dp.rf.rf[26][26] ),
    .X(_04045_));
 sky130_fd_sc_hd__o211ai_2 _09126_ (.A1(_01488_),
    .A2(\rvsingle.dp.rf.rf[27][26] ),
    .B1(_01491_),
    .C1(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__o211ai_2 _09127_ (.A1(_01106_),
    .A2(_04044_),
    .B1(_04046_),
    .C1(_01132_),
    .Y(_04047_));
 sky130_fd_sc_hd__o211ai_2 _09128_ (.A1(_01133_),
    .A2(_04042_),
    .B1(_04047_),
    .C1(_01117_),
    .Y(_04048_));
 sky130_fd_sc_hd__o311ai_2 _09129_ (.A1(_01117_),
    .A2(_04036_),
    .A3(_04041_),
    .B1(_01147_),
    .C1(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__nand4_2 _09130_ (.A(_01153_),
    .B(_04031_),
    .C(_04049_),
    .D(_01482_),
    .Y(_04050_));
 sky130_fd_sc_hd__o221a_2 _09131_ (.A1(_01066_),
    .A2(_01075_),
    .B1(_01482_),
    .B2(_01483_),
    .C1(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__a21oi_2 _09132_ (.A1(_01581_),
    .A2(_04050_),
    .B1(_01837_),
    .Y(_04052_));
 sky130_fd_sc_hd__nor4_2 _09133_ (.A(_04002_),
    .B(_04013_),
    .C(_04051_),
    .D(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__o22a_2 _09134_ (.A1(_04002_),
    .A2(_04013_),
    .B1(_04051_),
    .B2(_04052_),
    .X(_04054_));
 sky130_fd_sc_hd__or2_2 _09135_ (.A(_04053_),
    .B(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__nor2_2 _09136_ (.A(_03984_),
    .B(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__a21boi_2 _09137_ (.A1(_03909_),
    .A2(_03827_),
    .B1_N(_03908_),
    .Y(_04057_));
 sky130_fd_sc_hd__a221o_2 _09138_ (.A1(_03983_),
    .A2(_04053_),
    .B1(_04056_),
    .B2(_04057_),
    .C1(_03982_),
    .X(_04058_));
 sky130_fd_sc_hd__a31oi_2 _09139_ (.A1(_03775_),
    .A2(_03910_),
    .A3(_04056_),
    .B1(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__o22ai_2 _09140_ (.A1(_01348_),
    .A2(_01410_),
    .B1(_01415_),
    .B2(_04059_),
    .Y(_04060_));
 sky130_fd_sc_hd__a21o_2 _09141_ (.A1(_01182_),
    .A2(_01186_),
    .B1(_01249_),
    .X(_04061_));
 sky130_fd_sc_hd__and2_2 _09142_ (.A(_01250_),
    .B(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__nand2_2 _09143_ (.A(_04060_),
    .B(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__mux4_2 _09144_ (.A0(\rvsingle.dp.rf.rf[8][31] ),
    .A1(\rvsingle.dp.rf.rf[9][31] ),
    .A2(\rvsingle.dp.rf.rf[10][31] ),
    .A3(\rvsingle.dp.rf.rf[11][31] ),
    .S0(_01196_),
    .S1(_01203_),
    .X(_04064_));
 sky130_fd_sc_hd__or2_2 _09145_ (.A(_01196_),
    .B(\rvsingle.dp.rf.rf[12][31] ),
    .X(_04065_));
 sky130_fd_sc_hd__o211a_2 _09146_ (.A1(\rvsingle.dp.rf.rf[13][31] ),
    .A2(_01298_),
    .B1(_01311_),
    .C1(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__mux2_2 _09147_ (.A0(\rvsingle.dp.rf.rf[14][31] ),
    .A1(\rvsingle.dp.rf.rf[15][31] ),
    .S(_01196_),
    .X(_04067_));
 sky130_fd_sc_hd__a21o_2 _09148_ (.A1(_01226_),
    .A2(_04067_),
    .B1(_01210_),
    .X(_04068_));
 sky130_fd_sc_hd__o221a_2 _09149_ (.A1(_01232_),
    .A2(_04064_),
    .B1(_04066_),
    .B2(_04068_),
    .C1(_01224_),
    .X(_04069_));
 sky130_fd_sc_hd__mux4_2 _09150_ (.A0(\rvsingle.dp.rf.rf[4][31] ),
    .A1(\rvsingle.dp.rf.rf[5][31] ),
    .A2(\rvsingle.dp.rf.rf[6][31] ),
    .A3(\rvsingle.dp.rf.rf[7][31] ),
    .S0(_01225_),
    .S1(_01203_),
    .X(_04070_));
 sky130_fd_sc_hd__mux2_2 _09151_ (.A0(\rvsingle.dp.rf.rf[2][31] ),
    .A1(\rvsingle.dp.rf.rf[3][31] ),
    .S(_01196_),
    .X(_04071_));
 sky130_fd_sc_hd__or2_2 _09152_ (.A(_01195_),
    .B(\rvsingle.dp.rf.rf[0][31] ),
    .X(_04072_));
 sky130_fd_sc_hd__o211a_2 _09153_ (.A1(\rvsingle.dp.rf.rf[1][31] ),
    .A2(_01298_),
    .B1(_01311_),
    .C1(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__a211o_2 _09154_ (.A1(_01226_),
    .A2(_04071_),
    .B1(_04073_),
    .C1(_01232_),
    .X(_04074_));
 sky130_fd_sc_hd__o211a_2 _09155_ (.A1(_01210_),
    .A2(_04070_),
    .B1(_04074_),
    .C1(_01219_),
    .X(_04075_));
 sky130_fd_sc_hd__or3_2 _09156_ (.A(_01189_),
    .B(_04069_),
    .C(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__mux4_2 _09157_ (.A0(\rvsingle.dp.rf.rf[16][31] ),
    .A1(\rvsingle.dp.rf.rf[17][31] ),
    .A2(\rvsingle.dp.rf.rf[18][31] ),
    .A3(\rvsingle.dp.rf.rf[19][31] ),
    .S0(_01225_),
    .S1(_01226_),
    .X(_04077_));
 sky130_fd_sc_hd__mux4_2 _09158_ (.A0(\rvsingle.dp.rf.rf[20][31] ),
    .A1(\rvsingle.dp.rf.rf[21][31] ),
    .A2(\rvsingle.dp.rf.rf[22][31] ),
    .A3(\rvsingle.dp.rf.rf[23][31] ),
    .S0(_01225_),
    .S1(_01226_),
    .X(_04078_));
 sky130_fd_sc_hd__mux2_2 _09159_ (.A0(_04077_),
    .A1(_04078_),
    .S(_01232_),
    .X(_04079_));
 sky130_fd_sc_hd__or2_2 _09160_ (.A(_01225_),
    .B(\rvsingle.dp.rf.rf[28][31] ),
    .X(_04080_));
 sky130_fd_sc_hd__o211a_2 _09161_ (.A1(\rvsingle.dp.rf.rf[29][31] ),
    .A2(_01298_),
    .B1(_01311_),
    .C1(_04080_),
    .X(_04081_));
 sky130_fd_sc_hd__or2_2 _09162_ (.A(_01225_),
    .B(\rvsingle.dp.rf.rf[30][31] ),
    .X(_04082_));
 sky130_fd_sc_hd__o211a_2 _09163_ (.A1(_01298_),
    .A2(\rvsingle.dp.rf.rf[31][31] ),
    .B1(_01226_),
    .C1(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__mux4_2 _09164_ (.A0(\rvsingle.dp.rf.rf[24][31] ),
    .A1(\rvsingle.dp.rf.rf[25][31] ),
    .A2(\rvsingle.dp.rf.rf[26][31] ),
    .A3(\rvsingle.dp.rf.rf[27][31] ),
    .S0(_01196_),
    .S1(_01203_),
    .X(_04084_));
 sky130_fd_sc_hd__or2_2 _09165_ (.A(_01232_),
    .B(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__o311a_2 _09166_ (.A1(_01210_),
    .A2(_04081_),
    .A3(_04083_),
    .B1(_01224_),
    .C1(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__a211o_2 _09167_ (.A1(_01219_),
    .A2(_04079_),
    .B1(_01317_),
    .C1(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__mux4_2 _09168_ (.A0(\rvsingle.dp.rf.rf[24][31] ),
    .A1(\rvsingle.dp.rf.rf[25][31] ),
    .A2(\rvsingle.dp.rf.rf[26][31] ),
    .A3(\rvsingle.dp.rf.rf[27][31] ),
    .S0(_02212_),
    .S1(_01120_),
    .X(_04088_));
 sky130_fd_sc_hd__mux2_2 _09169_ (.A0(\rvsingle.dp.rf.rf[30][31] ),
    .A1(\rvsingle.dp.rf.rf[31][31] ),
    .S(_02212_),
    .X(_04089_));
 sky130_fd_sc_hd__or2_2 _09170_ (.A(_01100_),
    .B(\rvsingle.dp.rf.rf[28][31] ),
    .X(_04090_));
 sky130_fd_sc_hd__o211a_2 _09171_ (.A1(\rvsingle.dp.rf.rf[29][31] ),
    .A2(_01090_),
    .B1(_01094_),
    .C1(_04090_),
    .X(_04091_));
 sky130_fd_sc_hd__a211o_2 _09172_ (.A1(_01120_),
    .A2(_04089_),
    .B1(_01134_),
    .C1(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__o211a_2 _09173_ (.A1(_01114_),
    .A2(_04088_),
    .B1(_01118_),
    .C1(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__mux4_2 _09174_ (.A0(\rvsingle.dp.rf.rf[20][31] ),
    .A1(\rvsingle.dp.rf.rf[21][31] ),
    .A2(\rvsingle.dp.rf.rf[22][31] ),
    .A3(\rvsingle.dp.rf.rf[23][31] ),
    .S0(_02212_),
    .S1(_01120_),
    .X(_04094_));
 sky130_fd_sc_hd__or2_2 _09175_ (.A(_02212_),
    .B(\rvsingle.dp.rf.rf[18][31] ),
    .X(_04095_));
 sky130_fd_sc_hd__o211a_2 _09176_ (.A1(_01090_),
    .A2(\rvsingle.dp.rf.rf[19][31] ),
    .B1(_01120_),
    .C1(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__mux2_2 _09177_ (.A0(\rvsingle.dp.rf.rf[16][31] ),
    .A1(\rvsingle.dp.rf.rf[17][31] ),
    .S(_02212_),
    .X(_04097_));
 sky130_fd_sc_hd__a21o_2 _09178_ (.A1(_04097_),
    .A2(_01094_),
    .B1(_01114_),
    .X(_04098_));
 sky130_fd_sc_hd__o221a_2 _09179_ (.A1(_01134_),
    .A2(_04094_),
    .B1(_04096_),
    .B2(_04098_),
    .C1(_01157_),
    .X(_04099_));
 sky130_fd_sc_hd__mux4_2 _09180_ (.A0(\rvsingle.dp.rf.rf[12][31] ),
    .A1(\rvsingle.dp.rf.rf[13][31] ),
    .A2(\rvsingle.dp.rf.rf[14][31] ),
    .A3(\rvsingle.dp.rf.rf[15][31] ),
    .S0(_01100_),
    .S1(_01120_),
    .X(_04100_));
 sky130_fd_sc_hd__mux4_2 _09181_ (.A0(\rvsingle.dp.rf.rf[8][31] ),
    .A1(\rvsingle.dp.rf.rf[9][31] ),
    .A2(\rvsingle.dp.rf.rf[10][31] ),
    .A3(\rvsingle.dp.rf.rf[11][31] ),
    .S0(_01100_),
    .S1(_01120_),
    .X(_04101_));
 sky130_fd_sc_hd__mux2_2 _09182_ (.A0(_04100_),
    .A1(_04101_),
    .S(_01134_),
    .X(_04102_));
 sky130_fd_sc_hd__mux4_2 _09183_ (.A0(\rvsingle.dp.rf.rf[4][31] ),
    .A1(\rvsingle.dp.rf.rf[5][31] ),
    .A2(\rvsingle.dp.rf.rf[6][31] ),
    .A3(\rvsingle.dp.rf.rf[7][31] ),
    .S0(_02212_),
    .S1(_01120_),
    .X(_04103_));
 sky130_fd_sc_hd__mux2_2 _09184_ (.A0(\rvsingle.dp.rf.rf[2][31] ),
    .A1(\rvsingle.dp.rf.rf[3][31] ),
    .S(_01100_),
    .X(_04104_));
 sky130_fd_sc_hd__or2_2 _09185_ (.A(_01128_),
    .B(\rvsingle.dp.rf.rf[0][31] ),
    .X(_04105_));
 sky130_fd_sc_hd__o211a_2 _09186_ (.A1(\rvsingle.dp.rf.rf[1][31] ),
    .A2(_01090_),
    .B1(_01094_),
    .C1(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__a211o_2 _09187_ (.A1(_01120_),
    .A2(_04104_),
    .B1(_04106_),
    .C1(_01114_),
    .X(_04107_));
 sky130_fd_sc_hd__o211a_2 _09188_ (.A1(_01134_),
    .A2(_04103_),
    .B1(_04107_),
    .C1(_01157_),
    .X(_04108_));
 sky130_fd_sc_hd__a211o_2 _09189_ (.A1(_04102_),
    .A2(_01118_),
    .B1(_01147_),
    .C1(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__o311a_2 _09190_ (.A1(_01378_),
    .A2(_04093_),
    .A3(_04099_),
    .B1(_04109_),
    .C1(_01154_),
    .X(WriteData[31]));
 sky130_fd_sc_hd__a21o_2 _09191_ (.A1(_01085_),
    .A2(WriteData[31]),
    .B1(_01180_),
    .X(_04110_));
 sky130_fd_sc_hd__and4_2 _09192_ (.A(_01248_),
    .B(_04076_),
    .C(_04087_),
    .D(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__and3_2 _09193_ (.A(_01248_),
    .B(_04076_),
    .C(_04087_),
    .X(_04112_));
 sky130_fd_sc_hd__nor2_2 _09194_ (.A(_04112_),
    .B(_04110_),
    .Y(_04113_));
 sky130_fd_sc_hd__o21a_2 _09195_ (.A1(_04111_),
    .A2(_04113_),
    .B1(_01185_),
    .X(_04114_));
 sky130_fd_sc_hd__nor3_2 _09196_ (.A(_01185_),
    .B(_04111_),
    .C(_04113_),
    .Y(_04115_));
 sky130_fd_sc_hd__nor2_2 _09197_ (.A(_04114_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__or4b_2 _09198_ (.A(Instr[12]),
    .B(Instr[14]),
    .C(_01063_),
    .D_N(Instr[13]),
    .X(_04117_));
 sky130_fd_sc_hd__a31oi_2 _09199_ (.A1(_01250_),
    .A2(_04063_),
    .A3(_04116_),
    .B1(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__o2bb2ai_2 _09200_ (.A1_N(_01250_),
    .A2_N(_04063_),
    .B1(_04114_),
    .B2(_04115_),
    .Y(_04119_));
 sky130_fd_sc_hd__o21a_2 _09201_ (.A1(_02907_),
    .A2(_02963_),
    .B1(_02966_),
    .X(_04120_));
 sky130_fd_sc_hd__buf_1 _09202_ (.A(_01063_),
    .X(_04121_));
 sky130_fd_sc_hd__buf_1 _09203_ (.A(_01059_),
    .X(_04122_));
 sky130_fd_sc_hd__or2_2 _09204_ (.A(_04121_),
    .B(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__and3b_2 _09205_ (.A_N(_02962_),
    .B(_02964_),
    .C(_02965_),
    .X(_04124_));
 sky130_fd_sc_hd__o21ai_2 _09206_ (.A1(_01063_),
    .A2(_04122_),
    .B1(_04117_),
    .Y(_04125_));
 sky130_fd_sc_hd__nor2_2 _09207_ (.A(_02907_),
    .B(_02963_),
    .Y(_04126_));
 sky130_fd_sc_hd__o32a_2 _09208_ (.A1(_04121_),
    .A2(_04122_),
    .A3(_01066_),
    .B1(_04125_),
    .B2(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__o32a_2 _09209_ (.A1(_01060_),
    .A2(_04120_),
    .A3(_04123_),
    .B1(_04124_),
    .B2(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__inv_2 _09210_ (.A(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__a21oi_2 _09211_ (.A1(_04118_),
    .A2(_04119_),
    .B1(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_2 _09212_ (.A(_04110_),
    .B(_04112_),
    .Y(_04131_));
 sky130_fd_sc_hd__a211o_2 _09213_ (.A1(_04131_),
    .A2(_01066_),
    .B1(_04123_),
    .C1(_04113_),
    .X(_04132_));
 sky130_fd_sc_hd__a21boi_2 _09214_ (.A1(_04060_),
    .A2(_04062_),
    .B1_N(_01250_),
    .Y(_04133_));
 sky130_fd_sc_hd__nand3_2 _09215_ (.A(_01250_),
    .B(_04063_),
    .C(_04116_),
    .Y(_04134_));
 sky130_fd_sc_hd__o21a_2 _09216_ (.A1(_04121_),
    .A2(_04122_),
    .B1(_04117_),
    .X(_04135_));
 sky130_fd_sc_hd__buf_1 _09217_ (.A(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__buf_1 _09218_ (.A(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__o211ai_2 _09219_ (.A1(_04133_),
    .A2(_04116_),
    .B1(_04134_),
    .C1(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand3_2 _09220_ (.A(_04130_),
    .B(_04132_),
    .C(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__buf_1 _09221_ (.A(_02260_),
    .X(_04140_));
 sky130_fd_sc_hd__buf_1 _09222_ (.A(_01072_),
    .X(_04141_));
 sky130_fd_sc_hd__o2111a_2 _09223_ (.A1(_04140_),
    .A2(_04141_),
    .B1(Instr[13]),
    .C1(Instr[14]),
    .D1(_02259_),
    .X(_04142_));
 sky130_fd_sc_hd__buf_1 _09224_ (.A(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__o21ai_2 _09225_ (.A1(_01834_),
    .A2(_01838_),
    .B1(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__o41a_2 _09226_ (.A1(_01480_),
    .A2(_01453_),
    .A3(_01582_),
    .A4(_01579_),
    .B1(_01739_),
    .X(_04145_));
 sky130_fd_sc_hd__o21ba_2 _09227_ (.A1(_01740_),
    .A2(_01685_),
    .B1_N(_01737_),
    .X(_04146_));
 sky130_fd_sc_hd__or3b_2 _09228_ (.A(_04146_),
    .B(_01590_),
    .C_N(_01739_),
    .X(_04147_));
 sky130_fd_sc_hd__nor2_2 _09229_ (.A(_03231_),
    .B(_03406_),
    .Y(_04148_));
 sky130_fd_sc_hd__nor2_2 _09230_ (.A(_03573_),
    .B(_03735_),
    .Y(_04149_));
 sky130_fd_sc_hd__nand2_2 _09231_ (.A(_04148_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__a2bb2oi_2 _09232_ (.A1_N(_03047_),
    .A2_N(_03052_),
    .B1(_02967_),
    .B2(_03049_),
    .Y(_04151_));
 sky130_fd_sc_hd__o2111ai_2 _09233_ (.A1(_02851_),
    .A2(_02803_),
    .B1(_02856_),
    .C1(_02751_),
    .D1(_02861_),
    .Y(_04152_));
 sky130_fd_sc_hd__o2bb2ai_2 _09234_ (.A1_N(_02751_),
    .A2_N(_02857_),
    .B1(_04151_),
    .B2(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__o2111ai_2 _09235_ (.A1(_02374_),
    .A2(_02377_),
    .B1(_02464_),
    .C1(_02468_),
    .D1(_02475_),
    .Y(_04154_));
 sky130_fd_sc_hd__nand4_2 _09236_ (.A(_03056_),
    .B(_02576_),
    .C(_02661_),
    .D(_02667_),
    .Y(_04155_));
 sky130_fd_sc_hd__nor2_2 _09237_ (.A(_04154_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__a21o_2 _09238_ (.A1(_03056_),
    .A2(_02667_),
    .B1(_03057_),
    .X(_04157_));
 sky130_fd_sc_hd__o21bai_2 _09239_ (.A1(_04154_),
    .A2(_04157_),
    .B1_N(_03062_),
    .Y(_04158_));
 sky130_fd_sc_hd__a21oi_2 _09240_ (.A1(_04153_),
    .A2(_04156_),
    .B1(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__a21o_2 _09241_ (.A1(_03313_),
    .A2(_03405_),
    .B1(_03748_),
    .X(_04160_));
 sky130_fd_sc_hd__o21bai_2 _09242_ (.A1(_03231_),
    .A2(_04160_),
    .B1_N(_03753_),
    .Y(_04161_));
 sky130_fd_sc_hd__nand2_2 _09243_ (.A(_03572_),
    .B(_03755_),
    .Y(_04162_));
 sky130_fd_sc_hd__o21bai_2 _09244_ (.A1(_03735_),
    .A2(_04162_),
    .B1_N(_03756_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21oi_2 _09245_ (.A1(_04161_),
    .A2(_04149_),
    .B1(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__o21ai_2 _09246_ (.A1(_04150_),
    .A2(_04159_),
    .B1(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__and2_2 _09247_ (.A(_02184_),
    .B(_02265_),
    .X(_04166_));
 sky130_fd_sc_hd__a31oi_2 _09248_ (.A1(_04165_),
    .A2(_02101_),
    .A3(_04166_),
    .B1(_03768_),
    .Y(_04167_));
 sky130_fd_sc_hd__o22ai_2 _09249_ (.A1(_03770_),
    .A2(_04145_),
    .B1(_04147_),
    .B2(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__and2_2 _09250_ (.A(_01927_),
    .B(_01929_),
    .X(_04169_));
 sky130_fd_sc_hd__a21boi_2 _09251_ (.A1(_04168_),
    .A2(_04169_),
    .B1_N(_01927_),
    .Y(_04170_));
 sky130_fd_sc_hd__inv_2 _09252_ (.A(_01836_),
    .Y(_04171_));
 sky130_fd_sc_hd__nand2_2 _09253_ (.A(_04168_),
    .B(_04169_),
    .Y(_04172_));
 sky130_fd_sc_hd__o211ai_2 _09254_ (.A1(_04171_),
    .A2(_03772_),
    .B1(_01927_),
    .C1(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__o211ai_2 _09255_ (.A1(_01840_),
    .A2(_04170_),
    .B1(_04173_),
    .C1(_04137_),
    .Y(_04174_));
 sky130_fd_sc_hd__o21ai_2 _09256_ (.A1(_01804_),
    .A2(_04144_),
    .B1(_04174_),
    .Y(DataAdr[23]));
 sky130_fd_sc_hd__inv_2 _09257_ (.A(DataAdr[23]),
    .Y(_04175_));
 sky130_fd_sc_hd__nand3_2 _09258_ (.A(_03775_),
    .B(_03910_),
    .C(_04056_),
    .Y(_04176_));
 sky130_fd_sc_hd__a221oi_2 _09259_ (.A1(_03983_),
    .A2(_04053_),
    .B1(_04056_),
    .B2(_04057_),
    .C1(_03982_),
    .Y(_04177_));
 sky130_fd_sc_hd__a22oi_2 _09260_ (.A1(_01411_),
    .A2(_01412_),
    .B1(_04176_),
    .B2(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__o21bai_2 _09261_ (.A1(_01409_),
    .A2(_04178_),
    .B1_N(_01414_),
    .Y(_04179_));
 sky130_fd_sc_hd__and2_2 _09262_ (.A(_01411_),
    .B(_01412_),
    .X(_04180_));
 sky130_fd_sc_hd__o211ai_2 _09263_ (.A1(_04180_),
    .A2(_04059_),
    .B1(_01408_),
    .C1(_01414_),
    .Y(_04181_));
 sky130_fd_sc_hd__a21oi_2 _09264_ (.A1(_01185_),
    .A2(_01289_),
    .B1(_01347_),
    .Y(_04182_));
 sky130_fd_sc_hd__and4bb_2 _09265_ (.A_N(_04182_),
    .B_N(_04122_),
    .C(_04141_),
    .D(_01288_),
    .X(_04183_));
 sky130_fd_sc_hd__a31oi_2 _09266_ (.A1(_04179_),
    .A2(_04181_),
    .A3(_04137_),
    .B1(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__inv_2 _09267_ (.A(_04184_),
    .Y(DataAdr[29]));
 sky130_fd_sc_hd__nand2_2 _09268_ (.A(_01250_),
    .B(_04061_),
    .Y(_04185_));
 sky130_fd_sc_hd__o221ai_2 _09269_ (.A1(_01348_),
    .A2(_01410_),
    .B1(_01415_),
    .B2(_04059_),
    .C1(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__nand3_2 _09270_ (.A(_04063_),
    .B(_04137_),
    .C(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__a21oi_2 _09271_ (.A1(_01181_),
    .A2(_01185_),
    .B1(_01249_),
    .Y(_04188_));
 sky130_fd_sc_hd__or4b_2 _09272_ (.A(_04121_),
    .B(_04188_),
    .C(_04122_),
    .D_N(_01186_),
    .X(_04189_));
 sky130_fd_sc_hd__nand2_2 _09273_ (.A(_04187_),
    .B(_04189_),
    .Y(DataAdr[30]));
 sky130_fd_sc_hd__nor2_2 _09274_ (.A(DataAdr[29]),
    .B(DataAdr[30]),
    .Y(_04190_));
 sky130_fd_sc_hd__or2_2 _09275_ (.A(_04051_),
    .B(_04052_),
    .X(_04191_));
 sky130_fd_sc_hd__nand2_2 _09276_ (.A(_03909_),
    .B(_03827_),
    .Y(_04192_));
 sky130_fd_sc_hd__a22oi_2 _09277_ (.A1(_03908_),
    .A2(_04192_),
    .B1(_03775_),
    .B2(_03910_),
    .Y(_04193_));
 sky130_fd_sc_hd__o32ai_2 _09278_ (.A1(_04002_),
    .A2(_04013_),
    .A3(_04191_),
    .B1(_04055_),
    .B2(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hd__inv_2 _09279_ (.A(_03984_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_2 _09280_ (.A(_04194_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__inv_2 _09281_ (.A(_04053_),
    .Y(_04197_));
 sky130_fd_sc_hd__o211ai_2 _09282_ (.A1(_04055_),
    .A2(_04193_),
    .B1(_03984_),
    .C1(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__nand3_2 _09283_ (.A(_04196_),
    .B(_04198_),
    .C(_04137_),
    .Y(_04199_));
 sky130_fd_sc_hd__inv_2 _09284_ (.A(_03939_),
    .Y(_04200_));
 sky130_fd_sc_hd__o221ai_2 _09285_ (.A1(_01180_),
    .A2(_03978_),
    .B1(_03981_),
    .B2(_04200_),
    .C1(_04143_),
    .Y(_04201_));
 sky130_fd_sc_hd__o21ai_2 _09286_ (.A1(_04146_),
    .A2(_04167_),
    .B1(_01739_),
    .Y(_04202_));
 sky130_fd_sc_hd__nand3_2 _09287_ (.A(_01583_),
    .B(_01589_),
    .C(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__o211ai_2 _09288_ (.A1(_01742_),
    .A2(_04167_),
    .B1(_01590_),
    .C1(_01739_),
    .Y(_04204_));
 sky130_fd_sc_hd__o221a_2 _09289_ (.A1(_01585_),
    .A2(_01180_),
    .B1(_01586_),
    .B2(_01582_),
    .C1(_04143_),
    .X(_04205_));
 sky130_fd_sc_hd__a31oi_2 _09290_ (.A1(_04203_),
    .A2(_04204_),
    .A3(_04137_),
    .B1(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__nand3_2 _09291_ (.A(_04199_),
    .B(_04201_),
    .C(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__nor2_2 _09292_ (.A(_01925_),
    .B(_01928_),
    .Y(_04208_));
 sky130_fd_sc_hd__o211ai_2 _09293_ (.A1(_04169_),
    .A2(_04168_),
    .B1(_04137_),
    .C1(_04172_),
    .Y(_04209_));
 sky130_fd_sc_hd__o31a_2 _09294_ (.A1(_01898_),
    .A2(_04123_),
    .A3(_04208_),
    .B1(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__a21oi_2 _09295_ (.A1(_03741_),
    .A2(_02261_),
    .B1(_03727_),
    .Y(_04211_));
 sky130_fd_sc_hd__o21ai_2 _09296_ (.A1(_01737_),
    .A2(_01740_),
    .B1(_04143_),
    .Y(_04212_));
 sky130_fd_sc_hd__nand2_2 _09297_ (.A(_02015_),
    .B(_02016_),
    .Y(_04213_));
 sky130_fd_sc_hd__nand2_2 _09298_ (.A(_02098_),
    .B(_02100_),
    .Y(_04214_));
 sky130_fd_sc_hd__or3_2 _09299_ (.A(_04213_),
    .B(_04214_),
    .C(_03765_),
    .X(_04215_));
 sky130_fd_sc_hd__nand3_2 _09300_ (.A(_04165_),
    .B(_02101_),
    .C(_04166_),
    .Y(_04216_));
 sky130_fd_sc_hd__a31o_2 _09301_ (.A1(_04215_),
    .A2(_04216_),
    .A3(_03767_),
    .B1(_01742_),
    .X(_04217_));
 sky130_fd_sc_hd__a21oi_2 _09302_ (.A1(_04167_),
    .A2(_01742_),
    .B1(_04125_),
    .Y(_04218_));
 sky130_fd_sc_hd__a2bb2oi_2 _09303_ (.A1_N(_01685_),
    .A2_N(_04212_),
    .B1(_04217_),
    .B2(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__nand2_2 _09304_ (.A(_03648_),
    .B(_03650_),
    .Y(_04220_));
 sky130_fd_sc_hd__or2_2 _09305_ (.A(_03231_),
    .B(_03406_),
    .X(_04221_));
 sky130_fd_sc_hd__o21bai_2 _09306_ (.A1(_04221_),
    .A2(_04159_),
    .B1_N(_04161_),
    .Y(_04222_));
 sky130_fd_sc_hd__a22oi_2 _09307_ (.A1(_03572_),
    .A2(_03755_),
    .B1(_04222_),
    .B2(_03737_),
    .Y(_04223_));
 sky130_fd_sc_hd__o21ai_2 _09308_ (.A1(_04220_),
    .A2(_04223_),
    .B1(_03650_),
    .Y(_04224_));
 sky130_fd_sc_hd__nand2_2 _09309_ (.A(_04224_),
    .B(_03744_),
    .Y(_04225_));
 sky130_fd_sc_hd__nand2_2 _09310_ (.A(_03729_),
    .B(_03734_),
    .Y(_04226_));
 sky130_fd_sc_hd__o211ai_2 _09311_ (.A1(_04220_),
    .A2(_04223_),
    .B1(_04226_),
    .C1(_03650_),
    .Y(_04227_));
 sky130_fd_sc_hd__nand3_2 _09312_ (.A(_04225_),
    .B(_04136_),
    .C(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__o311a_2 _09313_ (.A1(_03731_),
    .A2(_04123_),
    .A3(_04211_),
    .B1(_04219_),
    .C1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__nor2_2 _09314_ (.A(_04002_),
    .B(_04013_),
    .Y(_04230_));
 sky130_fd_sc_hd__o21ai_2 _09315_ (.A1(_04230_),
    .A2(_04052_),
    .B1(_04143_),
    .Y(_04231_));
 sky130_fd_sc_hd__o21a_2 _09316_ (.A1(_04053_),
    .A2(_04054_),
    .B1(_04193_),
    .X(_04232_));
 sky130_fd_sc_hd__o21ai_2 _09317_ (.A1(_04055_),
    .A2(_04193_),
    .B1(_04136_),
    .Y(_04233_));
 sky130_fd_sc_hd__o22a_2 _09318_ (.A1(_04051_),
    .A2(_04231_),
    .B1(_04232_),
    .B2(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__nand3_2 _09319_ (.A(_04210_),
    .B(_04229_),
    .C(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__nor2_2 _09320_ (.A(_04207_),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__and4_2 _09321_ (.A(_01931_),
    .B(_02101_),
    .C(_02184_),
    .D(_02265_),
    .X(_04237_));
 sky130_fd_sc_hd__a21oi_2 _09322_ (.A1(_04165_),
    .A2(_04237_),
    .B1(_03774_),
    .Y(_04238_));
 sky130_fd_sc_hd__o21ai_2 _09323_ (.A1(_03830_),
    .A2(_04238_),
    .B1(_03827_),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2_2 _09324_ (.A(_03909_),
    .B(_03908_),
    .Y(_04240_));
 sky130_fd_sc_hd__inv_2 _09325_ (.A(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__nand2_2 _09326_ (.A(_04239_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__o211ai_2 _09327_ (.A1(_03830_),
    .A2(_04238_),
    .B1(_04240_),
    .C1(_03827_),
    .Y(_04243_));
 sky130_fd_sc_hd__a211o_2 _09328_ (.A1(_01581_),
    .A2(_03879_),
    .B1(_01066_),
    .C1(_01075_),
    .X(_04244_));
 sky130_fd_sc_hd__o31a_2 _09329_ (.A1(_01169_),
    .A2(_02259_),
    .A3(_01170_),
    .B1(_01063_),
    .X(_04245_));
 sky130_fd_sc_hd__or3b_2 _09330_ (.A(_04245_),
    .B(_04122_),
    .C_N(_02259_),
    .X(_04246_));
 sky130_fd_sc_hd__buf_1 _09331_ (.A(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__a211oi_2 _09332_ (.A1(_03907_),
    .A2(_04244_),
    .B1(_03881_),
    .C1(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__a31oi_2 _09333_ (.A1(_04242_),
    .A2(_04136_),
    .A3(_04243_),
    .B1(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__or3_2 _09334_ (.A(_02211_),
    .B(_02263_),
    .C(_03763_),
    .X(_04250_));
 sky130_fd_sc_hd__nand2_2 _09335_ (.A(_04165_),
    .B(_02265_),
    .Y(_04251_));
 sky130_fd_sc_hd__a21bo_2 _09336_ (.A1(_04250_),
    .A2(_04251_),
    .B1_N(_02184_),
    .X(_04252_));
 sky130_fd_sc_hd__nand3b_2 _09337_ (.A_N(_02184_),
    .B(_04250_),
    .C(_04251_),
    .Y(_04253_));
 sky130_fd_sc_hd__a31o_2 _09338_ (.A1(_01185_),
    .A2(_02261_),
    .A3(_02152_),
    .B1(_02181_),
    .X(_04254_));
 sky130_fd_sc_hd__and3_2 _09339_ (.A(_02151_),
    .B(_04254_),
    .C(_04143_),
    .X(_04255_));
 sky130_fd_sc_hd__a31oi_2 _09340_ (.A1(_04252_),
    .A2(_04253_),
    .A3(_04137_),
    .B1(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__inv_2 _09341_ (.A(_03565_),
    .Y(_04257_));
 sky130_fd_sc_hd__nand2_2 _09342_ (.A(_03565_),
    .B(_03567_),
    .Y(_04258_));
 sky130_fd_sc_hd__a21oi_2 _09343_ (.A1(_03064_),
    .A2(_04148_),
    .B1(_04161_),
    .Y(_04259_));
 sky130_fd_sc_hd__nor2_2 _09344_ (.A(_04258_),
    .B(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__o21a_2 _09345_ (.A1(_03454_),
    .A2(_03483_),
    .B1(_03572_),
    .X(_04261_));
 sky130_fd_sc_hd__o21ai_2 _09346_ (.A1(_04257_),
    .A2(_04260_),
    .B1(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__inv_2 _09347_ (.A(_04258_),
    .Y(_04263_));
 sky130_fd_sc_hd__a211o_2 _09348_ (.A1(_04222_),
    .A2(_04263_),
    .B1(_04257_),
    .C1(_04261_),
    .X(_04264_));
 sky130_fd_sc_hd__and3_2 _09349_ (.A(_01248_),
    .B(_03467_),
    .C(_03481_),
    .X(_04265_));
 sky130_fd_sc_hd__a2bb2o_2 _09350_ (.A1_N(_01066_),
    .A2_N(_01075_),
    .B1(_02261_),
    .B2(_03570_),
    .X(_04266_));
 sky130_fd_sc_hd__o211a_2 _09351_ (.A1(_04265_),
    .A2(_03454_),
    .B1(_04142_),
    .C1(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__a31oi_2 _09352_ (.A1(_04262_),
    .A2(_04264_),
    .A3(_04136_),
    .B1(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__a31oi_2 _09353_ (.A1(_01185_),
    .A2(_02261_),
    .A3(_03646_),
    .B1(_03649_),
    .Y(_04269_));
 sky130_fd_sc_hd__or3b_2 _09354_ (.A(_04121_),
    .B(_04122_),
    .C_N(_03645_),
    .X(_04270_));
 sky130_fd_sc_hd__o221ai_2 _09355_ (.A1(_03738_),
    .A2(_03739_),
    .B1(_03573_),
    .B2(_04259_),
    .C1(_04162_),
    .Y(_04271_));
 sky130_fd_sc_hd__o211ai_2 _09356_ (.A1(_04220_),
    .A2(_04223_),
    .B1(_04271_),
    .C1(_04136_),
    .Y(_04272_));
 sky130_fd_sc_hd__o21a_2 _09357_ (.A1(_04269_),
    .A2(_04270_),
    .B1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__nand4_2 _09358_ (.A(_04249_),
    .B(_04256_),
    .C(_04268_),
    .D(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__inv_2 _09359_ (.A(_02100_),
    .Y(_04275_));
 sky130_fd_sc_hd__nand3_2 _09360_ (.A(_04165_),
    .B(_02184_),
    .C(_02265_),
    .Y(_04276_));
 sky130_fd_sc_hd__a21oi_2 _09361_ (.A1(_03765_),
    .A2(_04276_),
    .B1(_04214_),
    .Y(_04277_));
 sky130_fd_sc_hd__o21bai_2 _09362_ (.A1(_04275_),
    .A2(_04277_),
    .B1_N(_04213_),
    .Y(_04278_));
 sky130_fd_sc_hd__inv_2 _09363_ (.A(_03765_),
    .Y(_04279_));
 sky130_fd_sc_hd__a31oi_2 _09364_ (.A1(_04165_),
    .A2(_02184_),
    .A3(_02265_),
    .B1(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__o211ai_2 _09365_ (.A1(_04214_),
    .A2(_04280_),
    .B1(_04213_),
    .C1(_02100_),
    .Y(_04281_));
 sky130_fd_sc_hd__a31oi_2 _09366_ (.A1(_01185_),
    .A2(_02261_),
    .A3(_02013_),
    .B1(_01959_),
    .Y(_04282_));
 sky130_fd_sc_hd__and4bb_2 _09367_ (.A_N(_04282_),
    .B_N(_04122_),
    .C(_04141_),
    .D(_02012_),
    .X(_04283_));
 sky130_fd_sc_hd__a31oi_2 _09368_ (.A1(_04278_),
    .A2(_04137_),
    .A3(_04281_),
    .B1(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__nor2_2 _09369_ (.A(_01185_),
    .B(_01405_),
    .Y(_04285_));
 sky130_fd_sc_hd__a211o_2 _09370_ (.A1(_01375_),
    .A2(_01406_),
    .B1(_04285_),
    .C1(_04247_),
    .X(_04286_));
 sky130_fd_sc_hd__nand2_2 _09371_ (.A(_04059_),
    .B(_04180_),
    .Y(_04287_));
 sky130_fd_sc_hd__o211ai_2 _09372_ (.A1(_04059_),
    .A2(_04180_),
    .B1(_04137_),
    .C1(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand3_2 _09373_ (.A(_04284_),
    .B(_04286_),
    .C(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__a31o_2 _09374_ (.A1(_04214_),
    .A2(_03765_),
    .A3(_04276_),
    .B1(_04125_),
    .X(_04290_));
 sky130_fd_sc_hd__o21a_2 _09375_ (.A1(_02081_),
    .A2(_02097_),
    .B1(_02068_),
    .X(_04291_));
 sky130_fd_sc_hd__a311o_2 _09376_ (.A1(_01837_),
    .A2(_01581_),
    .A3(_02067_),
    .B1(_04123_),
    .C1(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__o21ai_2 _09377_ (.A1(_04277_),
    .A2(_04290_),
    .B1(_04292_),
    .Y(DataAdr[18]));
 sky130_fd_sc_hd__inv_2 _09378_ (.A(DataAdr[18]),
    .Y(_04293_));
 sky130_fd_sc_hd__o21ai_2 _09379_ (.A1(_03143_),
    .A2(_03141_),
    .B1(_03230_),
    .Y(_04294_));
 sky130_fd_sc_hd__and2_2 _09380_ (.A(_03313_),
    .B(_03317_),
    .X(_04295_));
 sky130_fd_sc_hd__a41o_2 _09381_ (.A1(_03064_),
    .A2(_04295_),
    .A3(_03399_),
    .A4(_03405_),
    .B1(_03749_),
    .X(_04296_));
 sky130_fd_sc_hd__and2_2 _09382_ (.A(_03227_),
    .B(_03221_),
    .X(_04297_));
 sky130_fd_sc_hd__a21boi_2 _09383_ (.A1(_04296_),
    .A2(_04297_),
    .B1_N(_03227_),
    .Y(_04298_));
 sky130_fd_sc_hd__nand2_2 _09384_ (.A(_04296_),
    .B(_04297_),
    .Y(_04299_));
 sky130_fd_sc_hd__nand3_2 _09385_ (.A(_03227_),
    .B(_04294_),
    .C(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__o211ai_2 _09386_ (.A1(_04294_),
    .A2(_04298_),
    .B1(_04136_),
    .C1(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__o211ai_2 _09387_ (.A1(_03140_),
    .A2(_03143_),
    .B1(_04143_),
    .C1(_03112_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_2 _09388_ (.A(_03775_),
    .B(_03831_),
    .Y(_04303_));
 sky130_fd_sc_hd__a211o_2 _09389_ (.A1(_04165_),
    .A2(_04237_),
    .B1(_03774_),
    .C1(_03831_),
    .X(_04304_));
 sky130_fd_sc_hd__nand3_2 _09390_ (.A(_04303_),
    .B(_04304_),
    .C(_04136_),
    .Y(_04305_));
 sky130_fd_sc_hd__o211ai_2 _09391_ (.A1(_03825_),
    .A2(_03803_),
    .B1(_04143_),
    .C1(_03826_),
    .Y(_04306_));
 sky130_fd_sc_hd__and4_2 _09392_ (.A(_04301_),
    .B(_04302_),
    .C(_04305_),
    .D(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__o21ai_2 _09393_ (.A1(_04155_),
    .A2(_03054_),
    .B1(_04157_),
    .Y(_04308_));
 sky130_fd_sc_hd__and2_2 _09394_ (.A(_02464_),
    .B(_02475_),
    .X(_04309_));
 sky130_fd_sc_hd__nand2_2 _09395_ (.A(_04308_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__o21ai_2 _09396_ (.A1(_02377_),
    .A2(_02374_),
    .B1(_02468_),
    .Y(_04311_));
 sky130_fd_sc_hd__a21oi_2 _09397_ (.A1(_02464_),
    .A2(_04310_),
    .B1(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__a31o_2 _09398_ (.A1(_04311_),
    .A2(_02464_),
    .A3(_04310_),
    .B1(_04125_),
    .X(_04313_));
 sky130_fd_sc_hd__o21a_2 _09399_ (.A1(_02317_),
    .A2(_02377_),
    .B1(_02373_),
    .X(_04314_));
 sky130_fd_sc_hd__a2bb2o_2 _09400_ (.A1_N(_04312_),
    .A2_N(_04313_),
    .B1(_04314_),
    .B2(_04143_),
    .X(DataAdr[7]));
 sky130_fd_sc_hd__o21a_2 _09401_ (.A1(_04297_),
    .A2(_04296_),
    .B1(_04135_),
    .X(_04315_));
 sky130_fd_sc_hd__o211a_2 _09402_ (.A1(_03222_),
    .A2(_03220_),
    .B1(_04142_),
    .C1(_03223_),
    .X(_04316_));
 sky130_fd_sc_hd__a21o_2 _09403_ (.A1(_04315_),
    .A2(_04299_),
    .B1(_04316_),
    .X(DataAdr[10]));
 sky130_fd_sc_hd__nor2_2 _09404_ (.A(DataAdr[7]),
    .B(DataAdr[10]),
    .Y(_04317_));
 sky130_fd_sc_hd__o21ai_2 _09405_ (.A1(_04263_),
    .A2(_04222_),
    .B1(_04135_),
    .Y(_04318_));
 sky130_fd_sc_hd__and3_2 _09406_ (.A(_03561_),
    .B(_01185_),
    .C(_02261_),
    .X(_04319_));
 sky130_fd_sc_hd__and3_2 _09407_ (.A(Instr[13]),
    .B(Instr[14]),
    .C(_04141_),
    .X(_04320_));
 sky130_fd_sc_hd__o211ai_2 _09408_ (.A1(_03513_),
    .A2(_04319_),
    .B1(_03564_),
    .C1(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__o21ai_2 _09409_ (.A1(_04260_),
    .A2(_04318_),
    .B1(_04321_),
    .Y(DataAdr[12]));
 sky130_fd_sc_hd__a211o_2 _09410_ (.A1(_02257_),
    .A2(_01085_),
    .B1(_01837_),
    .C1(_03142_),
    .X(_04322_));
 sky130_fd_sc_hd__a21o_2 _09411_ (.A1(_02211_),
    .A2(_04322_),
    .B1(_04247_),
    .X(_04323_));
 sky130_fd_sc_hd__o2111ai_2 _09412_ (.A1(_02265_),
    .A2(_04165_),
    .B1(_04247_),
    .C1(_04117_),
    .D1(_04251_),
    .Y(_04324_));
 sky130_fd_sc_hd__o21ai_2 _09413_ (.A1(_02263_),
    .A2(_04323_),
    .B1(_04324_),
    .Y(DataAdr[16]));
 sky130_fd_sc_hd__nand2_2 _09414_ (.A(_03064_),
    .B(_04295_),
    .Y(_04325_));
 sky130_fd_sc_hd__nand2_2 _09415_ (.A(_03399_),
    .B(_03405_),
    .Y(_04326_));
 sky130_fd_sc_hd__a21oi_2 _09416_ (.A1(_03313_),
    .A2(_04325_),
    .B1(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__a31o_2 _09417_ (.A1(_03313_),
    .A2(_04326_),
    .A3(_04325_),
    .B1(_04125_),
    .X(_04328_));
 sky130_fd_sc_hd__a211o_2 _09418_ (.A1(_03398_),
    .A2(_03402_),
    .B1(_04247_),
    .C1(_03366_),
    .X(_04329_));
 sky130_fd_sc_hd__o21ai_2 _09419_ (.A1(_04327_),
    .A2(_04328_),
    .B1(_04329_),
    .Y(DataAdr[9]));
 sky130_fd_sc_hd__a221o_2 _09420_ (.A1(_03313_),
    .A2(_03317_),
    .B1(_04153_),
    .B2(_04156_),
    .C1(_04158_),
    .X(_04330_));
 sky130_fd_sc_hd__o211a_2 _09421_ (.A1(_03311_),
    .A2(_03316_),
    .B1(_04142_),
    .C1(_03312_),
    .X(_04331_));
 sky130_fd_sc_hd__a31o_2 _09422_ (.A1(_04325_),
    .A2(_04330_),
    .A3(_04135_),
    .B1(_04331_),
    .X(DataAdr[8]));
 sky130_fd_sc_hd__o21ai_2 _09423_ (.A1(_02854_),
    .A2(_02750_),
    .B1(_02855_),
    .Y(_04332_));
 sky130_fd_sc_hd__and2_2 _09424_ (.A(_02751_),
    .B(_02856_),
    .X(_04333_));
 sky130_fd_sc_hd__o21ai_2 _09425_ (.A1(_02803_),
    .A2(_02851_),
    .B1(_02861_),
    .Y(_04334_));
 sky130_fd_sc_hd__o22ai_2 _09426_ (.A1(_02803_),
    .A2(_02851_),
    .B1(_04334_),
    .B2(_04151_),
    .Y(_04335_));
 sky130_fd_sc_hd__o21ai_2 _09427_ (.A1(_04333_),
    .A2(_04335_),
    .B1(_04135_),
    .Y(_04336_));
 sky130_fd_sc_hd__and3_2 _09428_ (.A(_02751_),
    .B(_02856_),
    .C(_04335_),
    .X(_04337_));
 sky130_fd_sc_hd__o22ai_2 _09429_ (.A1(_04247_),
    .A2(_04332_),
    .B1(_04336_),
    .B2(_04337_),
    .Y(DataAdr[3]));
 sky130_fd_sc_hd__o21ai_2 _09430_ (.A1(_03047_),
    .A2(_03052_),
    .B1(_03049_),
    .Y(_04338_));
 sky130_fd_sc_hd__o211a_2 _09431_ (.A1(_03047_),
    .A2(_03052_),
    .B1(_02967_),
    .C1(_03049_),
    .X(_04339_));
 sky130_fd_sc_hd__a211o_2 _09432_ (.A1(_04120_),
    .A2(_04338_),
    .B1(_04125_),
    .C1(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__or2_2 _09433_ (.A(_04334_),
    .B(_04151_),
    .X(_04341_));
 sky130_fd_sc_hd__a21oi_2 _09434_ (.A1(_04151_),
    .A2(_04334_),
    .B1(_04125_),
    .Y(_04342_));
 sky130_fd_sc_hd__o211a_2 _09435_ (.A1(_02848_),
    .A2(_02803_),
    .B1(_02850_),
    .C1(_04142_),
    .X(_04343_));
 sky130_fd_sc_hd__a21oi_2 _09436_ (.A1(_04341_),
    .A2(_04342_),
    .B1(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__nand4_2 _09437_ (.A(_04340_),
    .B(_04344_),
    .C(_01069_),
    .D(_01067_),
    .Y(_04345_));
 sky130_fd_sc_hd__a221o_2 _09438_ (.A1(_02751_),
    .A2(_02857_),
    .B1(_02862_),
    .B2(_03053_),
    .C1(_02577_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_2 _09439_ (.A(_04153_),
    .B(_02577_),
    .Y(_04347_));
 sky130_fd_sc_hd__o211a_2 _09440_ (.A1(_02570_),
    .A2(_02534_),
    .B1(_02572_),
    .C1(_04142_),
    .X(_04348_));
 sky130_fd_sc_hd__a31o_2 _09441_ (.A1(_04346_),
    .A2(_04135_),
    .A3(_04347_),
    .B1(_04348_),
    .X(DataAdr[4]));
 sky130_fd_sc_hd__nor3_2 _09442_ (.A(DataAdr[3]),
    .B(_04345_),
    .C(DataAdr[4]),
    .Y(_04349_));
 sky130_fd_sc_hd__nand2_2 _09443_ (.A(_02661_),
    .B(_02667_),
    .Y(_04350_));
 sky130_fd_sc_hd__a21o_2 _09444_ (.A1(_03056_),
    .A2(_04347_),
    .B1(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__o211ai_2 _09445_ (.A1(_02534_),
    .A2(_02573_),
    .B1(_04350_),
    .C1(_04347_),
    .Y(_04352_));
 sky130_fd_sc_hd__o211a_2 _09446_ (.A1(_02665_),
    .A2(_02660_),
    .B1(_04320_),
    .C1(_02666_),
    .X(_04353_));
 sky130_fd_sc_hd__a31oi_2 _09447_ (.A1(_04351_),
    .A2(_04136_),
    .A3(_04352_),
    .B1(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__and3_2 _09448_ (.A(_03056_),
    .B(_02576_),
    .C(_02667_),
    .X(_04355_));
 sky130_fd_sc_hd__a311o_2 _09449_ (.A1(_04153_),
    .A2(_02661_),
    .A3(_04355_),
    .B1(_03058_),
    .C1(_04309_),
    .X(_04356_));
 sky130_fd_sc_hd__o211a_2 _09450_ (.A1(_02463_),
    .A2(_02472_),
    .B1(_02432_),
    .C1(_04142_),
    .X(_04357_));
 sky130_fd_sc_hd__a31oi_2 _09451_ (.A1(_04310_),
    .A2(_04356_),
    .A3(_04136_),
    .B1(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__nand4b_2 _09452_ (.A_N(DataAdr[8]),
    .B(_04349_),
    .C(_04354_),
    .D(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__nor4_2 _09453_ (.A(DataAdr[12]),
    .B(DataAdr[16]),
    .C(DataAdr[9]),
    .D(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand4_2 _09454_ (.A(_04293_),
    .B(_04307_),
    .C(_04317_),
    .D(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__nor3_2 _09455_ (.A(_04274_),
    .B(_04289_),
    .C(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__nand4_2 _09456_ (.A(_04175_),
    .B(_04190_),
    .C(_04236_),
    .D(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__buf_1 _09457_ (.A(_04140_),
    .X(_04364_));
 sky130_fd_sc_hd__buf_1 _09458_ (.A(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__o21bai_2 _09459_ (.A1(_04139_),
    .A2(_04363_),
    .B1_N(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__buf_1 _09460_ (.A(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__nand2_2 _09461_ (.A(_02914_),
    .B(_02913_),
    .Y(_04368_));
 sky130_fd_sc_hd__o21ai_2 _09462_ (.A1(_04140_),
    .A2(_01069_),
    .B1(_01067_),
    .Y(_04369_));
 sky130_fd_sc_hd__and3_2 _09463_ (.A(_04368_),
    .B(PC[0]),
    .C(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__nand2_2 _09464_ (.A(PC[1]),
    .B(_03045_),
    .Y(_04371_));
 sky130_fd_sc_hd__o211ai_2 _09465_ (.A1(_01094_),
    .A2(_01069_),
    .B1(_03044_),
    .C1(_01058_),
    .Y(_04372_));
 sky130_fd_sc_hd__and2_2 _09466_ (.A(_04371_),
    .B(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__o21ai_2 _09467_ (.A1(_04370_),
    .A2(_04373_),
    .B1(_04366_),
    .Y(_04374_));
 sky130_fd_sc_hd__o21ai_2 _09468_ (.A1(_01058_),
    .A2(_04367_),
    .B1(_04374_),
    .Y(_00622_));
 sky130_fd_sc_hd__buf_1 _09469_ (.A(PC[0]),
    .X(_04375_));
 sky130_fd_sc_hd__buf_1 _09470_ (.A(_04375_),
    .X(_00621_));
 sky130_fd_sc_hd__and4b_2 _09471_ (.A_N(_01067_),
    .B(_02912_),
    .C(_01071_),
    .D(_01062_),
    .X(_04376_));
 sky130_fd_sc_hd__buf_1 _09472_ (.A(_04376_),
    .X(MemWrite));
 sky130_fd_sc_hd__buf_1 _09473_ (.A(_01154_),
    .X(_04377_));
 sky130_fd_sc_hd__and3_2 _09474_ (.A(_04377_),
    .B(_02885_),
    .C(_02906_),
    .X(_04378_));
 sky130_fd_sc_hd__buf_1 _09475_ (.A(_04378_),
    .X(WriteData[0]));
 sky130_fd_sc_hd__and3_2 _09476_ (.A(_01154_),
    .B(_03956_),
    .C(_03977_),
    .X(_04379_));
 sky130_fd_sc_hd__buf_1 _09477_ (.A(_04379_),
    .X(WriteData[27]));
 sky130_fd_sc_hd__o211ai_2 _09478_ (.A1(_01962_),
    .A2(_02212_),
    .B1(_04049_),
    .C1(_04031_),
    .Y(_04380_));
 sky130_fd_sc_hd__inv_2 _09479_ (.A(_04380_),
    .Y(WriteData[26]));
 sky130_fd_sc_hd__and3_2 _09480_ (.A(_01154_),
    .B(_03790_),
    .C(_03801_),
    .X(_04381_));
 sky130_fd_sc_hd__buf_1 _09481_ (.A(_04381_),
    .X(WriteData[24]));
 sky130_fd_sc_hd__and3_2 _09482_ (.A(_01154_),
    .B(_01774_),
    .C(_01802_),
    .X(_04382_));
 sky130_fd_sc_hd__buf_1 _09483_ (.A(_04382_),
    .X(WriteData[23]));
 sky130_fd_sc_hd__and3_2 _09484_ (.A(_01154_),
    .B(_01869_),
    .C(_01896_),
    .X(_04383_));
 sky130_fd_sc_hd__buf_1 _09485_ (.A(_04383_),
    .X(WriteData[22]));
 sky130_fd_sc_hd__and3_2 _09486_ (.A(_04377_),
    .B(_01536_),
    .C(_01577_),
    .X(_04384_));
 sky130_fd_sc_hd__buf_1 _09487_ (.A(_04384_),
    .X(WriteData[21]));
 sky130_fd_sc_hd__and3_2 _09488_ (.A(_01154_),
    .B(_01641_),
    .C(_01683_),
    .X(_04385_));
 sky130_fd_sc_hd__buf_1 _09489_ (.A(_04385_),
    .X(WriteData[20]));
 sky130_fd_sc_hd__inv_2 _09490_ (.A(_02011_),
    .Y(WriteData[19]));
 sky130_fd_sc_hd__inv_2 _09491_ (.A(_02065_),
    .Y(WriteData[18]));
 sky130_fd_sc_hd__inv_2 _09492_ (.A(_02150_),
    .Y(WriteData[17]));
 sky130_fd_sc_hd__inv_2 _09493_ (.A(_02257_),
    .Y(WriteData[16]));
 sky130_fd_sc_hd__inv_2 _09494_ (.A(_03697_),
    .Y(WriteData[15]));
 sky130_fd_sc_hd__inv_2 _09495_ (.A(_03644_),
    .Y(WriteData[14]));
 sky130_fd_sc_hd__inv_2 _09496_ (.A(_03453_),
    .Y(WriteData[13]));
 sky130_fd_sc_hd__and3_2 _09497_ (.A(_04377_),
    .B(_03537_),
    .C(_03560_),
    .X(_04386_));
 sky130_fd_sc_hd__buf_1 _09498_ (.A(_04386_),
    .X(WriteData[12]));
 sky130_fd_sc_hd__inv_2 _09499_ (.A(_03111_),
    .Y(WriteData[11]));
 sky130_fd_sc_hd__and3_2 _09500_ (.A(_04377_),
    .B(_03194_),
    .C(_03217_),
    .X(_04387_));
 sky130_fd_sc_hd__buf_1 _09501_ (.A(_04387_),
    .X(WriteData[10]));
 sky130_fd_sc_hd__and3_2 _09502_ (.A(_04377_),
    .B(_03341_),
    .C(_03364_),
    .X(_04388_));
 sky130_fd_sc_hd__buf_1 _09503_ (.A(_04388_),
    .X(WriteData[9]));
 sky130_fd_sc_hd__o211ai_2 _09504_ (.A1(_01962_),
    .A2(_02212_),
    .B1(_03280_),
    .C1(_03255_),
    .Y(_04389_));
 sky130_fd_sc_hd__inv_2 _09505_ (.A(_04389_),
    .Y(WriteData[8]));
 sky130_fd_sc_hd__and3_2 _09506_ (.A(_04377_),
    .B(_02346_),
    .C(_02371_),
    .X(_04390_));
 sky130_fd_sc_hd__buf_1 _09507_ (.A(_04390_),
    .X(WriteData[7]));
 sky130_fd_sc_hd__inv_2 _09508_ (.A(_02427_),
    .Y(WriteData[6]));
 sky130_fd_sc_hd__inv_2 _09509_ (.A(_02662_),
    .Y(WriteData[5]));
 sky130_fd_sc_hd__and3_2 _09510_ (.A(_04377_),
    .B(_02504_),
    .C(_02529_),
    .X(_04391_));
 sky130_fd_sc_hd__buf_1 _09511_ (.A(_04391_),
    .X(WriteData[4]));
 sky130_fd_sc_hd__and3_2 _09512_ (.A(_04377_),
    .B(_02721_),
    .C(_02745_),
    .X(_04392_));
 sky130_fd_sc_hd__buf_1 _09513_ (.A(_04392_),
    .X(WriteData[3]));
 sky130_fd_sc_hd__and3_2 _09514_ (.A(_04377_),
    .B(_02774_),
    .C(_02797_),
    .X(_04393_));
 sky130_fd_sc_hd__buf_1 _09515_ (.A(_04393_),
    .X(WriteData[2]));
 sky130_fd_sc_hd__and3_2 _09516_ (.A(_04377_),
    .B(_03019_),
    .C(_03042_),
    .X(_04394_));
 sky130_fd_sc_hd__buf_1 _09517_ (.A(_04394_),
    .X(WriteData[1]));
 sky130_fd_sc_hd__inv_2 _09518_ (.A(_04130_),
    .Y(DataAdr[0]));
 sky130_fd_sc_hd__o211ai_2 _09519_ (.A1(_03050_),
    .A2(_03047_),
    .B1(_03051_),
    .C1(_04143_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand2_2 _09520_ (.A(_04340_),
    .B(_04395_),
    .Y(DataAdr[1]));
 sky130_fd_sc_hd__inv_2 _09521_ (.A(_04344_),
    .Y(DataAdr[2]));
 sky130_fd_sc_hd__inv_2 _09522_ (.A(_04354_),
    .Y(DataAdr[5]));
 sky130_fd_sc_hd__inv_2 _09523_ (.A(_04358_),
    .Y(DataAdr[6]));
 sky130_fd_sc_hd__nand2_2 _09524_ (.A(_04301_),
    .B(_04302_),
    .Y(DataAdr[11]));
 sky130_fd_sc_hd__inv_2 _09525_ (.A(_04268_),
    .Y(DataAdr[13]));
 sky130_fd_sc_hd__inv_2 _09526_ (.A(_04273_),
    .Y(DataAdr[14]));
 sky130_fd_sc_hd__or4_2 _09527_ (.A(_04121_),
    .B(_04122_),
    .C(_03731_),
    .D(_04211_),
    .X(_04396_));
 sky130_fd_sc_hd__nand2_2 _09528_ (.A(_04228_),
    .B(_04396_),
    .Y(DataAdr[15]));
 sky130_fd_sc_hd__inv_2 _09529_ (.A(_04256_),
    .Y(DataAdr[17]));
 sky130_fd_sc_hd__inv_2 _09530_ (.A(_04284_),
    .Y(DataAdr[19]));
 sky130_fd_sc_hd__inv_2 _09531_ (.A(_04219_),
    .Y(DataAdr[20]));
 sky130_fd_sc_hd__inv_2 _09532_ (.A(_04206_),
    .Y(DataAdr[21]));
 sky130_fd_sc_hd__inv_2 _09533_ (.A(_04210_),
    .Y(DataAdr[22]));
 sky130_fd_sc_hd__nand2_2 _09534_ (.A(_04305_),
    .B(_04306_),
    .Y(DataAdr[24]));
 sky130_fd_sc_hd__inv_2 _09535_ (.A(_04249_),
    .Y(DataAdr[25]));
 sky130_fd_sc_hd__inv_2 _09536_ (.A(_04234_),
    .Y(DataAdr[26]));
 sky130_fd_sc_hd__nand2_2 _09537_ (.A(_04199_),
    .B(_04201_),
    .Y(DataAdr[27]));
 sky130_fd_sc_hd__nand2_2 _09538_ (.A(_04288_),
    .B(_04286_),
    .Y(DataAdr[28]));
 sky130_fd_sc_hd__nand2_2 _09539_ (.A(_04138_),
    .B(_04132_),
    .Y(DataAdr[31]));
 sky130_fd_sc_hd__buf_1 _09540_ (.A(PC[2]),
    .X(_04397_));
 sky130_fd_sc_hd__buf_1 _09541_ (.A(_04366_),
    .X(_04398_));
 sky130_fd_sc_hd__nand4_2 _09542_ (.A(_04368_),
    .B(PC[0]),
    .C(_04369_),
    .D(_04372_),
    .Y(_04399_));
 sky130_fd_sc_hd__nand2_2 _09543_ (.A(_04371_),
    .B(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__o211a_2 _09544_ (.A1(_01114_),
    .A2(_01069_),
    .B1(_04397_),
    .C1(_02800_),
    .X(_04401_));
 sky130_fd_sc_hd__nor2_2 _09545_ (.A(_04397_),
    .B(_02801_),
    .Y(_04402_));
 sky130_fd_sc_hd__or2_2 _09546_ (.A(_04401_),
    .B(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__xnor2_2 _09547_ (.A(_04400_),
    .B(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2_2 _09548_ (.A(_04398_),
    .B(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__o21ai_2 _09549_ (.A1(_04397_),
    .A2(_04367_),
    .B1(_04405_),
    .Y(\rvsingle.dp.PCNext[2] ));
 sky130_fd_sc_hd__xnor2_2 _09550_ (.A(_04397_),
    .B(PC[3]),
    .Y(_04406_));
 sky130_fd_sc_hd__nor2_2 _09551_ (.A(PC[3]),
    .B(_02748_),
    .Y(_04407_));
 sky130_fd_sc_hd__nand2_2 _09552_ (.A(PC[3]),
    .B(_02748_),
    .Y(_04408_));
 sky130_fd_sc_hd__and2b_2 _09553_ (.A_N(_04407_),
    .B(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__a2bb2oi_2 _09554_ (.A1_N(_04397_),
    .A2_N(_02801_),
    .B1(_04371_),
    .B2(_04399_),
    .Y(_04410_));
 sky130_fd_sc_hd__a21o_2 _09555_ (.A1(_04397_),
    .A2(_02801_),
    .B1(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__xor2_2 _09556_ (.A(_04409_),
    .B(_04411_),
    .X(_04412_));
 sky130_fd_sc_hd__nand2_2 _09557_ (.A(_04398_),
    .B(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__o21ai_2 _09558_ (.A1(_04367_),
    .A2(_04406_),
    .B1(_04413_),
    .Y(\rvsingle.dp.PCNext[3] ));
 sky130_fd_sc_hd__o211a_2 _09559_ (.A1(Instr[11]),
    .A2(_01078_),
    .B1(PC[4]),
    .C1(_02531_),
    .X(_04414_));
 sky130_fd_sc_hd__nor2_2 _09560_ (.A(PC[4]),
    .B(_02532_),
    .Y(_04415_));
 sky130_fd_sc_hd__or2_2 _09561_ (.A(_04414_),
    .B(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__o22ai_2 _09562_ (.A1(PC[3]),
    .A2(_02748_),
    .B1(_04401_),
    .B2(_04410_),
    .Y(_04417_));
 sky130_fd_sc_hd__and3_2 _09563_ (.A(_04408_),
    .B(_04416_),
    .C(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__a21oi_2 _09564_ (.A1(_04408_),
    .A2(_04417_),
    .B1(_04416_),
    .Y(_04419_));
 sky130_fd_sc_hd__nor2_2 _09565_ (.A(_04418_),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__and3_2 _09566_ (.A(PC[2]),
    .B(PC[3]),
    .C(PC[4]),
    .X(_04421_));
 sky130_fd_sc_hd__buf_1 _09567_ (.A(_04139_),
    .X(_04422_));
 sky130_fd_sc_hd__buf_1 _09568_ (.A(_04363_),
    .X(_04423_));
 sky130_fd_sc_hd__a21o_2 _09569_ (.A1(_04397_),
    .A2(PC[3]),
    .B1(PC[4]),
    .X(_04424_));
 sky130_fd_sc_hd__buf_1 _09570_ (.A(_01080_),
    .X(_04425_));
 sky130_fd_sc_hd__buf_1 _09571_ (.A(_04425_),
    .X(_04426_));
 sky130_fd_sc_hd__buf_1 _09572_ (.A(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__o211ai_2 _09573_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04424_),
    .C1(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__o2bb2ai_2 _09574_ (.A1_N(_04367_),
    .A2_N(_04420_),
    .B1(_04421_),
    .B2(_04428_),
    .Y(\rvsingle.dp.PCNext[4] ));
 sky130_fd_sc_hd__buf_1 _09575_ (.A(PC[5]),
    .X(_04429_));
 sky130_fd_sc_hd__nand2_2 _09576_ (.A(_04429_),
    .B(_04421_),
    .Y(_04430_));
 sky130_fd_sc_hd__a31o_2 _09577_ (.A1(_04397_),
    .A2(PC[3]),
    .A3(PC[4]),
    .B1(_04429_),
    .X(_04431_));
 sky130_fd_sc_hd__nand2_2 _09578_ (.A(_04430_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__or2_2 _09579_ (.A(Instr[25]),
    .B(_04429_),
    .X(_04433_));
 sky130_fd_sc_hd__nand2_2 _09580_ (.A(Instr[25]),
    .B(_04429_),
    .Y(_04434_));
 sky130_fd_sc_hd__o211ai_2 _09581_ (.A1(_04414_),
    .A2(_04419_),
    .B1(_04433_),
    .C1(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__a221o_2 _09582_ (.A1(PC[4]),
    .A2(_02532_),
    .B1(_04433_),
    .B2(_04434_),
    .C1(_04419_),
    .X(_04436_));
 sky130_fd_sc_hd__nand3_2 _09583_ (.A(_04366_),
    .B(_04435_),
    .C(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__o21ai_2 _09584_ (.A1(_04367_),
    .A2(_04432_),
    .B1(_04437_),
    .Y(\rvsingle.dp.PCNext[5] ));
 sky130_fd_sc_hd__xor2_2 _09585_ (.A(Instr[26]),
    .B(PC[6]),
    .X(_04438_));
 sky130_fd_sc_hd__a22o_2 _09586_ (.A1(Instr[25]),
    .A2(_04429_),
    .B1(_02532_),
    .B2(PC[4]),
    .X(_04439_));
 sky130_fd_sc_hd__o22a_2 _09587_ (.A1(Instr[25]),
    .A2(_04429_),
    .B1(_04439_),
    .B2(_04419_),
    .X(_04440_));
 sky130_fd_sc_hd__nor2_2 _09588_ (.A(_04438_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__o221a_2 _09589_ (.A1(Instr[25]),
    .A2(_04429_),
    .B1(_04439_),
    .B2(_04419_),
    .C1(_04438_),
    .X(_04442_));
 sky130_fd_sc_hd__nor2_2 _09590_ (.A(_04441_),
    .B(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__and3_2 _09591_ (.A(_04429_),
    .B(PC[6]),
    .C(_04421_),
    .X(_04444_));
 sky130_fd_sc_hd__a41o_2 _09592_ (.A1(_04397_),
    .A2(PC[3]),
    .A3(PC[4]),
    .A4(_04429_),
    .B1(PC[6]),
    .X(_04445_));
 sky130_fd_sc_hd__o211ai_2 _09593_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04445_),
    .C1(_04427_),
    .Y(_04446_));
 sky130_fd_sc_hd__o2bb2ai_2 _09594_ (.A1_N(_04367_),
    .A2_N(_04443_),
    .B1(_04444_),
    .B2(_04446_),
    .Y(\rvsingle.dp.PCNext[6] ));
 sky130_fd_sc_hd__nand2_2 _09595_ (.A(Instr[27]),
    .B(PC[7]),
    .Y(_04447_));
 sky130_fd_sc_hd__or2_2 _09596_ (.A(Instr[27]),
    .B(PC[7]),
    .X(_04448_));
 sky130_fd_sc_hd__nand2_2 _09597_ (.A(_04447_),
    .B(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__a21oi_2 _09598_ (.A1(Instr[26]),
    .A2(PC[6]),
    .B1(_04442_),
    .Y(_04450_));
 sky130_fd_sc_hd__xnor2_2 _09599_ (.A(_04449_),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__o21a_2 _09600_ (.A1(_04139_),
    .A2(_04363_),
    .B1(_04426_),
    .X(_04452_));
 sky130_fd_sc_hd__buf_1 _09601_ (.A(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__buf_1 _09602_ (.A(_04139_),
    .X(_04454_));
 sky130_fd_sc_hd__buf_1 _09603_ (.A(_04363_),
    .X(_04455_));
 sky130_fd_sc_hd__and4_2 _09604_ (.A(PC[5]),
    .B(PC[6]),
    .C(PC[7]),
    .D(_04421_),
    .X(_04456_));
 sky130_fd_sc_hd__nor2_2 _09605_ (.A(PC[7]),
    .B(_04444_),
    .Y(_04457_));
 sky130_fd_sc_hd__nor2_2 _09606_ (.A(_04456_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__buf_1 _09607_ (.A(_04427_),
    .X(_04459_));
 sky130_fd_sc_hd__o211ai_2 _09608_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04458_),
    .C1(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__o21ai_2 _09609_ (.A1(_04451_),
    .A2(_04453_),
    .B1(_04460_),
    .Y(\rvsingle.dp.PCNext[7] ));
 sky130_fd_sc_hd__and3_2 _09610_ (.A(_04438_),
    .B(_04447_),
    .C(_04448_),
    .X(_04461_));
 sky130_fd_sc_hd__o221ai_2 _09611_ (.A1(Instr[25]),
    .A2(_04429_),
    .B1(_04439_),
    .B2(_04419_),
    .C1(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__and3_2 _09612_ (.A(_04448_),
    .B(PC[6]),
    .C(Instr[26]),
    .X(_04463_));
 sky130_fd_sc_hd__a21oi_2 _09613_ (.A1(Instr[27]),
    .A2(PC[7]),
    .B1(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__and2_2 _09614_ (.A(_04462_),
    .B(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__xnor2_2 _09615_ (.A(Instr[28]),
    .B(PC[8]),
    .Y(_04466_));
 sky130_fd_sc_hd__xnor2_2 _09616_ (.A(_04465_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__xor2_2 _09617_ (.A(PC[8]),
    .B(_04456_),
    .X(_04468_));
 sky130_fd_sc_hd__o211ai_2 _09618_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04468_),
    .C1(_04459_),
    .Y(_04469_));
 sky130_fd_sc_hd__o21ai_2 _09619_ (.A1(_04467_),
    .A2(_04453_),
    .B1(_04469_),
    .Y(\rvsingle.dp.PCNext[8] ));
 sky130_fd_sc_hd__and2_2 _09620_ (.A(Instr[29]),
    .B(PC[9]),
    .X(_04470_));
 sky130_fd_sc_hd__nor2_2 _09621_ (.A(Instr[29]),
    .B(PC[9]),
    .Y(_04471_));
 sky130_fd_sc_hd__nor2_2 _09622_ (.A(_04470_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__o2bb2a_2 _09623_ (.A1_N(Instr[28]),
    .A2_N(PC[8]),
    .B1(_04465_),
    .B2(_04466_),
    .X(_04473_));
 sky130_fd_sc_hd__xor2_2 _09624_ (.A(_04472_),
    .B(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__and3_2 _09625_ (.A(PC[8]),
    .B(PC[9]),
    .C(_04456_),
    .X(_04475_));
 sky130_fd_sc_hd__a21oi_2 _09626_ (.A1(PC[8]),
    .A2(_04456_),
    .B1(PC[9]),
    .Y(_04476_));
 sky130_fd_sc_hd__nor2_2 _09627_ (.A(_04475_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__o211ai_2 _09628_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04477_),
    .C1(_04459_),
    .Y(_04478_));
 sky130_fd_sc_hd__o21ai_2 _09629_ (.A1(_04474_),
    .A2(_04453_),
    .B1(_04478_),
    .Y(\rvsingle.dp.PCNext[9] ));
 sky130_fd_sc_hd__xor2_2 _09630_ (.A(PC[10]),
    .B(_04475_),
    .X(_04479_));
 sky130_fd_sc_hd__inv_2 _09631_ (.A(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__nand2_2 _09632_ (.A(Instr[30]),
    .B(PC[10]),
    .Y(_04481_));
 sky130_fd_sc_hd__or2_2 _09633_ (.A(Instr[30]),
    .B(PC[10]),
    .X(_04482_));
 sky130_fd_sc_hd__or2_2 _09634_ (.A(Instr[29]),
    .B(PC[9]),
    .X(_04483_));
 sky130_fd_sc_hd__a31o_2 _09635_ (.A1(_04483_),
    .A2(PC[8]),
    .A3(Instr[28]),
    .B1(_04470_),
    .X(_04484_));
 sky130_fd_sc_hd__or3_2 _09636_ (.A(_04470_),
    .B(_04471_),
    .C(_04466_),
    .X(_04485_));
 sky130_fd_sc_hd__a21oi_2 _09637_ (.A1(_04462_),
    .A2(_04464_),
    .B1(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__a211o_2 _09638_ (.A1(_04481_),
    .A2(_04482_),
    .B1(_04484_),
    .C1(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__nand2_2 _09639_ (.A(_04481_),
    .B(_04482_),
    .Y(_04488_));
 sky130_fd_sc_hd__o21bai_2 _09640_ (.A1(_04484_),
    .A2(_04486_),
    .B1_N(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__nand3_2 _09641_ (.A(_04366_),
    .B(_04487_),
    .C(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__o21ai_2 _09642_ (.A1(_04367_),
    .A2(_04480_),
    .B1(_04490_),
    .Y(\rvsingle.dp.PCNext[10] ));
 sky130_fd_sc_hd__o21ai_2 _09643_ (.A1(_04140_),
    .A2(MemWrite),
    .B1(_01090_),
    .Y(_04491_));
 sky130_fd_sc_hd__o31a_2 _09644_ (.A1(Instr[7]),
    .A2(_04140_),
    .A3(MemWrite),
    .B1(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__mux2_2 _09645_ (.A0(_04492_),
    .A1(Instr[31]),
    .S(_04369_),
    .X(_04493_));
 sky130_fd_sc_hd__and2_2 _09646_ (.A(PC[11]),
    .B(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__nor2_2 _09647_ (.A(PC[11]),
    .B(_04493_),
    .Y(_04495_));
 sky130_fd_sc_hd__or2_2 _09648_ (.A(_04494_),
    .B(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__a21oi_2 _09649_ (.A1(_04481_),
    .A2(_04489_),
    .B1(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__and3_2 _09650_ (.A(_04481_),
    .B(_04489_),
    .C(_04496_),
    .X(_04498_));
 sky130_fd_sc_hd__or2_2 _09651_ (.A(_04497_),
    .B(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__and3_2 _09652_ (.A(PC[10]),
    .B(PC[11]),
    .C(_04475_),
    .X(_04500_));
 sky130_fd_sc_hd__a21oi_2 _09653_ (.A1(PC[10]),
    .A2(_04475_),
    .B1(PC[11]),
    .Y(_04501_));
 sky130_fd_sc_hd__nor2_2 _09654_ (.A(_04500_),
    .B(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__o211ai_2 _09655_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04502_),
    .C1(_04459_),
    .Y(_04503_));
 sky130_fd_sc_hd__o21ai_2 _09656_ (.A1(_04499_),
    .A2(_04453_),
    .B1(_04503_),
    .Y(\rvsingle.dp.PCNext[11] ));
 sky130_fd_sc_hd__a21oi_2 _09657_ (.A1(PC[11]),
    .A2(_04493_),
    .B1(_04497_),
    .Y(_04504_));
 sky130_fd_sc_hd__buf_1 _09658_ (.A(_02912_),
    .X(_04505_));
 sky130_fd_sc_hd__buf_1 _09659_ (.A(_01175_),
    .X(_04506_));
 sky130_fd_sc_hd__buf_1 _09660_ (.A(_01171_),
    .X(_04507_));
 sky130_fd_sc_hd__a31o_2 _09661_ (.A1(Instr[12]),
    .A2(_04505_),
    .A3(_04506_),
    .B1(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__and2_2 _09662_ (.A(_04508_),
    .B(PC[12]),
    .X(_04509_));
 sky130_fd_sc_hd__nor2_2 _09663_ (.A(PC[12]),
    .B(_04508_),
    .Y(_04510_));
 sky130_fd_sc_hd__or2_2 _09664_ (.A(_04509_),
    .B(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__xnor2_2 _09665_ (.A(_04504_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__xor2_2 _09666_ (.A(PC[12]),
    .B(_04500_),
    .X(_04513_));
 sky130_fd_sc_hd__o211ai_2 _09667_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04513_),
    .C1(_04459_),
    .Y(_04514_));
 sky130_fd_sc_hd__o21ai_2 _09668_ (.A1(_04512_),
    .A2(_04453_),
    .B1(_04514_),
    .Y(\rvsingle.dp.PCNext[12] ));
 sky130_fd_sc_hd__and3_2 _09669_ (.A(Instr[13]),
    .B(_02912_),
    .C(_04506_),
    .X(_04515_));
 sky130_fd_sc_hd__o21a_2 _09670_ (.A1(_04507_),
    .A2(_04515_),
    .B1(PC[13]),
    .X(_04516_));
 sky130_fd_sc_hd__a311o_2 _09671_ (.A1(Instr[13]),
    .A2(_02912_),
    .A3(_04506_),
    .B1(_04507_),
    .C1(PC[13]),
    .X(_04517_));
 sky130_fd_sc_hd__or2b_2 _09672_ (.A(_04516_),
    .B_N(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__o21ba_2 _09673_ (.A1(_04511_),
    .A2(_04504_),
    .B1_N(_04509_),
    .X(_04519_));
 sky130_fd_sc_hd__xnor2_2 _09674_ (.A(_04518_),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__and3_2 _09675_ (.A(PC[12]),
    .B(PC[13]),
    .C(_04500_),
    .X(_04521_));
 sky130_fd_sc_hd__buf_1 _09676_ (.A(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__a21oi_2 _09677_ (.A1(PC[12]),
    .A2(_04500_),
    .B1(PC[13]),
    .Y(_04523_));
 sky130_fd_sc_hd__nor2_2 _09678_ (.A(_04522_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__o211ai_2 _09679_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04524_),
    .C1(_04459_),
    .Y(_04525_));
 sky130_fd_sc_hd__o21ai_2 _09680_ (.A1(_04520_),
    .A2(_04453_),
    .B1(_04525_),
    .Y(\rvsingle.dp.PCNext[13] ));
 sky130_fd_sc_hd__or3_2 _09681_ (.A(_04509_),
    .B(_04510_),
    .C(_04518_),
    .X(_04526_));
 sky130_fd_sc_hd__o21bai_2 _09682_ (.A1(_04494_),
    .A2(_04497_),
    .B1_N(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__a21oi_2 _09683_ (.A1(_04509_),
    .A2(_04517_),
    .B1(_04516_),
    .Y(_04528_));
 sky130_fd_sc_hd__a31o_2 _09684_ (.A1(Instr[14]),
    .A2(_04505_),
    .A3(_04506_),
    .B1(_04507_),
    .X(_04529_));
 sky130_fd_sc_hd__xnor2_2 _09685_ (.A(PC[14]),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__a21oi_2 _09686_ (.A1(_04527_),
    .A2(_04528_),
    .B1(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__o311a_2 _09687_ (.A1(_04511_),
    .A2(_04518_),
    .A3(_04504_),
    .B1(_04528_),
    .C1(_04530_),
    .X(_04532_));
 sky130_fd_sc_hd__or2_2 _09688_ (.A(_04531_),
    .B(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__xor2_2 _09689_ (.A(PC[14]),
    .B(_04522_),
    .X(_04534_));
 sky130_fd_sc_hd__o211ai_2 _09690_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04534_),
    .C1(_04459_),
    .Y(_04535_));
 sky130_fd_sc_hd__o21ai_2 _09691_ (.A1(_04533_),
    .A2(_04453_),
    .B1(_04535_),
    .Y(\rvsingle.dp.PCNext[14] ));
 sky130_fd_sc_hd__a31o_2 _09692_ (.A1(_01225_),
    .A2(_04505_),
    .A3(_04506_),
    .B1(_04507_),
    .X(_04536_));
 sky130_fd_sc_hd__nand2_2 _09693_ (.A(_04536_),
    .B(PC[15]),
    .Y(_04537_));
 sky130_fd_sc_hd__a311o_2 _09694_ (.A1(_01225_),
    .A2(_04505_),
    .A3(_04506_),
    .B1(_04507_),
    .C1(PC[15]),
    .X(_04538_));
 sky130_fd_sc_hd__nand2_2 _09695_ (.A(_04537_),
    .B(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__a21oi_2 _09696_ (.A1(PC[14]),
    .A2(_04529_),
    .B1(_04531_),
    .Y(_04540_));
 sky130_fd_sc_hd__xnor2_2 _09697_ (.A(_04539_),
    .B(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a21oi_2 _09698_ (.A1(PC[14]),
    .A2(_04522_),
    .B1(PC[15]),
    .Y(_04542_));
 sky130_fd_sc_hd__and3_2 _09699_ (.A(PC[14]),
    .B(PC[15]),
    .C(_04522_),
    .X(_04543_));
 sky130_fd_sc_hd__nor2_2 _09700_ (.A(_04542_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__o211ai_2 _09701_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04544_),
    .C1(_04459_),
    .Y(_04545_));
 sky130_fd_sc_hd__o21ai_2 _09702_ (.A1(_04541_),
    .A2(_04453_),
    .B1(_04545_),
    .Y(\rvsingle.dp.PCNext[15] ));
 sky130_fd_sc_hd__a31o_2 _09703_ (.A1(_01226_),
    .A2(_02912_),
    .A3(_01175_),
    .B1(_01171_),
    .X(_04546_));
 sky130_fd_sc_hd__xnor2_2 _09704_ (.A(PC[16]),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__and3_2 _09705_ (.A(_04538_),
    .B(PC[14]),
    .C(_04529_),
    .X(_04548_));
 sky130_fd_sc_hd__a21o_2 _09706_ (.A1(PC[15]),
    .A2(_04536_),
    .B1(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__or2_2 _09707_ (.A(_04530_),
    .B(_04539_),
    .X(_04550_));
 sky130_fd_sc_hd__a21oi_2 _09708_ (.A1(_04527_),
    .A2(_04528_),
    .B1(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hd__nor2_2 _09709_ (.A(_04549_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__xnor2_2 _09710_ (.A(_04547_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__and4_2 _09711_ (.A(PC[14]),
    .B(PC[15]),
    .C(PC[16]),
    .D(_04522_),
    .X(_04554_));
 sky130_fd_sc_hd__nor2_2 _09712_ (.A(PC[16]),
    .B(_04543_),
    .Y(_04555_));
 sky130_fd_sc_hd__nor2_2 _09713_ (.A(_04554_),
    .B(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__o211ai_2 _09714_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04556_),
    .C1(_04459_),
    .Y(_04557_));
 sky130_fd_sc_hd__o21ai_2 _09715_ (.A1(_04553_),
    .A2(_04453_),
    .B1(_04557_),
    .Y(\rvsingle.dp.PCNext[16] ));
 sky130_fd_sc_hd__o21a_2 _09716_ (.A1(_04507_),
    .A2(_01176_),
    .B1(PC[17]),
    .X(_04558_));
 sky130_fd_sc_hd__a311o_2 _09717_ (.A1(_01232_),
    .A2(_02912_),
    .A3(_01175_),
    .B1(_01171_),
    .C1(PC[17]),
    .X(_04559_));
 sky130_fd_sc_hd__or2b_2 _09718_ (.A(_04558_),
    .B_N(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__nor2_2 _09719_ (.A(_04547_),
    .B(_04552_),
    .Y(_04561_));
 sky130_fd_sc_hd__a21oi_2 _09720_ (.A1(PC[16]),
    .A2(_04546_),
    .B1(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__xnor2_2 _09721_ (.A(_04560_),
    .B(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__nand2_2 _09722_ (.A(PC[17]),
    .B(_04554_),
    .Y(_04564_));
 sky130_fd_sc_hd__a41o_2 _09723_ (.A1(PC[14]),
    .A2(PC[15]),
    .A3(PC[16]),
    .A4(_04522_),
    .B1(PC[17]),
    .X(_04565_));
 sky130_fd_sc_hd__nand2_2 _09724_ (.A(_04564_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__o211a_2 _09725_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04566_),
    .C1(_04427_),
    .X(_04567_));
 sky130_fd_sc_hd__a21oi_2 _09726_ (.A1(_04398_),
    .A2(_04563_),
    .B1(_04567_),
    .Y(\rvsingle.dp.PCNext[17] ));
 sky130_fd_sc_hd__a31o_2 _09727_ (.A1(_04559_),
    .A2(PC[16]),
    .A3(_04546_),
    .B1(_04558_),
    .X(_04568_));
 sky130_fd_sc_hd__a21oi_2 _09728_ (.A1(_04561_),
    .A2(_04559_),
    .B1(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__a31o_2 _09729_ (.A1(_01224_),
    .A2(_02912_),
    .A3(_01175_),
    .B1(_04507_),
    .X(_04570_));
 sky130_fd_sc_hd__nand2_2 _09730_ (.A(_04570_),
    .B(PC[18]),
    .Y(_04571_));
 sky130_fd_sc_hd__a311o_2 _09731_ (.A1(_01224_),
    .A2(_02912_),
    .A3(_04506_),
    .B1(_04507_),
    .C1(PC[18]),
    .X(_04572_));
 sky130_fd_sc_hd__nand2_2 _09732_ (.A(_04571_),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__xnor2_2 _09733_ (.A(_04569_),
    .B(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__xnor2_2 _09734_ (.A(PC[18]),
    .B(_04564_),
    .Y(_04575_));
 sky130_fd_sc_hd__o211ai_2 _09735_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04575_),
    .C1(_04459_),
    .Y(_04576_));
 sky130_fd_sc_hd__o21ai_2 _09736_ (.A1(_04574_),
    .A2(_04453_),
    .B1(_04576_),
    .Y(\rvsingle.dp.PCNext[18] ));
 sky130_fd_sc_hd__a31o_2 _09737_ (.A1(_01189_),
    .A2(_02912_),
    .A3(_01175_),
    .B1(_04507_),
    .X(_04577_));
 sky130_fd_sc_hd__xnor2_2 _09738_ (.A(PC[19]),
    .B(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__o21ai_2 _09739_ (.A1(_04573_),
    .A2(_04569_),
    .B1(_04571_),
    .Y(_04579_));
 sky130_fd_sc_hd__xor2_2 _09740_ (.A(_04578_),
    .B(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__a31oi_2 _09741_ (.A1(PC[17]),
    .A2(PC[18]),
    .A3(_04554_),
    .B1(PC[19]),
    .Y(_04581_));
 sky130_fd_sc_hd__and4_2 _09742_ (.A(PC[17]),
    .B(PC[18]),
    .C(PC[19]),
    .D(_04554_),
    .X(_04582_));
 sky130_fd_sc_hd__or2_2 _09743_ (.A(_04581_),
    .B(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__o211a_2 _09744_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04583_),
    .C1(_04427_),
    .X(_04584_));
 sky130_fd_sc_hd__a21oi_2 _09745_ (.A1(_04398_),
    .A2(_04580_),
    .B1(_04584_),
    .Y(\rvsingle.dp.PCNext[19] ));
 sky130_fd_sc_hd__or4_2 _09746_ (.A(_04547_),
    .B(_04560_),
    .C(_04573_),
    .D(_04578_),
    .X(_04585_));
 sky130_fd_sc_hd__a22o_2 _09747_ (.A1(_04577_),
    .A2(PC[19]),
    .B1(PC[18]),
    .B2(_04570_),
    .X(_04586_));
 sky130_fd_sc_hd__a21o_2 _09748_ (.A1(_04568_),
    .A2(_04572_),
    .B1(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__o21ai_2 _09749_ (.A1(PC[19]),
    .A2(_04577_),
    .B1(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__o21ai_2 _09750_ (.A1(_04585_),
    .A2(_04552_),
    .B1(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__buf_1 _09751_ (.A(Instr[31]),
    .X(_04590_));
 sky130_fd_sc_hd__and2_2 _09752_ (.A(_04590_),
    .B(PC[20]),
    .X(_04591_));
 sky130_fd_sc_hd__or2_2 _09753_ (.A(Instr[31]),
    .B(PC[20]),
    .X(_04592_));
 sky130_fd_sc_hd__or2b_2 _09754_ (.A(_04591_),
    .B_N(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__xor2_2 _09755_ (.A(_04589_),
    .B(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__xor2_2 _09756_ (.A(PC[20]),
    .B(_04582_),
    .X(_04595_));
 sky130_fd_sc_hd__o211ai_2 _09757_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04595_),
    .C1(_04427_),
    .Y(_04596_));
 sky130_fd_sc_hd__o21ai_2 _09758_ (.A1(_04594_),
    .A2(_04452_),
    .B1(_04596_),
    .Y(\rvsingle.dp.PCNext[20] ));
 sky130_fd_sc_hd__and3_2 _09759_ (.A(PC[20]),
    .B(PC[21]),
    .C(_04582_),
    .X(_04597_));
 sky130_fd_sc_hd__a21oi_2 _09760_ (.A1(PC[20]),
    .A2(_04582_),
    .B1(PC[21]),
    .Y(_04598_));
 sky130_fd_sc_hd__or2_2 _09761_ (.A(_04597_),
    .B(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__xnor2_2 _09762_ (.A(Instr[31]),
    .B(PC[21]),
    .Y(_04600_));
 sky130_fd_sc_hd__a21oi_2 _09763_ (.A1(_04589_),
    .A2(_04592_),
    .B1(_04591_),
    .Y(_04601_));
 sky130_fd_sc_hd__xor2_2 _09764_ (.A(_04600_),
    .B(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__nand2_2 _09765_ (.A(_04398_),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__o21ai_2 _09766_ (.A1(_04367_),
    .A2(_04599_),
    .B1(_04603_),
    .Y(\rvsingle.dp.PCNext[21] ));
 sky130_fd_sc_hd__nor2_2 _09767_ (.A(_04593_),
    .B(_04600_),
    .Y(_04604_));
 sky130_fd_sc_hd__o21a_2 _09768_ (.A1(PC[20]),
    .A2(PC[21]),
    .B1(_04590_),
    .X(_04605_));
 sky130_fd_sc_hd__a21oi_2 _09769_ (.A1(_04589_),
    .A2(_04604_),
    .B1(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__and2_2 _09770_ (.A(_04590_),
    .B(PC[22]),
    .X(_04607_));
 sky130_fd_sc_hd__nor2_2 _09771_ (.A(_04590_),
    .B(PC[22]),
    .Y(_04608_));
 sky130_fd_sc_hd__or2_2 _09772_ (.A(_04607_),
    .B(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__xnor2_2 _09773_ (.A(_04606_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__and4_2 _09774_ (.A(PC[20]),
    .B(PC[21]),
    .C(PC[22]),
    .D(_04582_),
    .X(_04611_));
 sky130_fd_sc_hd__buf_1 _09775_ (.A(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__nor2_2 _09776_ (.A(PC[22]),
    .B(_04597_),
    .Y(_04613_));
 sky130_fd_sc_hd__nor2_2 _09777_ (.A(_04612_),
    .B(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__o211ai_2 _09778_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04614_),
    .C1(_04427_),
    .Y(_04615_));
 sky130_fd_sc_hd__o21ai_2 _09779_ (.A1(_04610_),
    .A2(_04452_),
    .B1(_04615_),
    .Y(\rvsingle.dp.PCNext[22] ));
 sky130_fd_sc_hd__xnor2_2 _09780_ (.A(PC[23]),
    .B(_04612_),
    .Y(_04616_));
 sky130_fd_sc_hd__buf_1 _09781_ (.A(_04590_),
    .X(_04617_));
 sky130_fd_sc_hd__buf_1 _09782_ (.A(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__nand2_2 _09783_ (.A(_04590_),
    .B(PC[23]),
    .Y(_04619_));
 sky130_fd_sc_hd__or2_2 _09784_ (.A(_04590_),
    .B(PC[23]),
    .X(_04620_));
 sky130_fd_sc_hd__nor2_2 _09785_ (.A(_04609_),
    .B(_04606_),
    .Y(_04621_));
 sky130_fd_sc_hd__a221o_2 _09786_ (.A1(_04618_),
    .A2(PC[22]),
    .B1(_04619_),
    .B2(_04620_),
    .C1(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__o211ai_2 _09787_ (.A1(_04607_),
    .A2(_04621_),
    .B1(_04619_),
    .C1(_04620_),
    .Y(_04623_));
 sky130_fd_sc_hd__nand3_2 _09788_ (.A(_04366_),
    .B(_04622_),
    .C(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__o21ai_2 _09789_ (.A1(_04398_),
    .A2(_04616_),
    .B1(_04624_),
    .Y(\rvsingle.dp.PCNext[23] ));
 sky130_fd_sc_hd__or3b_2 _09790_ (.A(_04591_),
    .B(_04600_),
    .C_N(_04592_),
    .X(_04625_));
 sky130_fd_sc_hd__nand2_2 _09791_ (.A(_04619_),
    .B(_04620_),
    .Y(_04626_));
 sky130_fd_sc_hd__or4_2 _09792_ (.A(_04585_),
    .B(_04625_),
    .C(_04609_),
    .D(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__o21bai_2 _09793_ (.A1(_04549_),
    .A2(_04551_),
    .B1_N(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__or4_2 _09794_ (.A(_04588_),
    .B(_04625_),
    .C(_04609_),
    .D(_04626_),
    .X(_04629_));
 sky130_fd_sc_hd__or4bb_2 _09795_ (.A(_04605_),
    .B(_04607_),
    .C_N(_04619_),
    .D_N(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__inv_2 _09796_ (.A(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__nand2_2 _09797_ (.A(_04617_),
    .B(PC[24]),
    .Y(_04632_));
 sky130_fd_sc_hd__or2_2 _09798_ (.A(_04590_),
    .B(PC[24]),
    .X(_04633_));
 sky130_fd_sc_hd__nand2_2 _09799_ (.A(_04632_),
    .B(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__a21o_2 _09800_ (.A1(_04628_),
    .A2(_04631_),
    .B1(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__o21ai_2 _09801_ (.A1(_04627_),
    .A2(_04552_),
    .B1(_04631_),
    .Y(_04636_));
 sky130_fd_sc_hd__a21o_2 _09802_ (.A1(_04632_),
    .A2(_04633_),
    .B1(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__nand2_2 _09803_ (.A(_04635_),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__and3_2 _09804_ (.A(PC[23]),
    .B(PC[24]),
    .C(_04612_),
    .X(_04639_));
 sky130_fd_sc_hd__a21oi_2 _09805_ (.A1(PC[23]),
    .A2(_04612_),
    .B1(PC[24]),
    .Y(_04640_));
 sky130_fd_sc_hd__nor2_2 _09806_ (.A(_04639_),
    .B(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__o211ai_2 _09807_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04641_),
    .C1(_04427_),
    .Y(_04642_));
 sky130_fd_sc_hd__o21ai_2 _09808_ (.A1(_04638_),
    .A2(_04452_),
    .B1(_04642_),
    .Y(\rvsingle.dp.PCNext[24] ));
 sky130_fd_sc_hd__xnor2_2 _09809_ (.A(PC[25]),
    .B(_04639_),
    .Y(_04643_));
 sky130_fd_sc_hd__xnor2_2 _09810_ (.A(_04617_),
    .B(PC[25]),
    .Y(_04644_));
 sky130_fd_sc_hd__nand3_2 _09811_ (.A(_04632_),
    .B(_04635_),
    .C(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__a21o_2 _09812_ (.A1(_04632_),
    .A2(_04635_),
    .B1(_04644_),
    .X(_04646_));
 sky130_fd_sc_hd__nand3_2 _09813_ (.A(_04366_),
    .B(_04645_),
    .C(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__o21ai_2 _09814_ (.A1(_04398_),
    .A2(_04643_),
    .B1(_04647_),
    .Y(\rvsingle.dp.PCNext[25] ));
 sky130_fd_sc_hd__nor2_2 _09815_ (.A(_04644_),
    .B(_04634_),
    .Y(_04648_));
 sky130_fd_sc_hd__o21a_2 _09816_ (.A1(PC[24]),
    .A2(PC[25]),
    .B1(_04617_),
    .X(_04649_));
 sky130_fd_sc_hd__a21oi_2 _09817_ (.A1(_04636_),
    .A2(_04648_),
    .B1(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__nand2_2 _09818_ (.A(_04590_),
    .B(PC[26]),
    .Y(_04651_));
 sky130_fd_sc_hd__or2_2 _09819_ (.A(_04590_),
    .B(PC[26]),
    .X(_04652_));
 sky130_fd_sc_hd__nand2_2 _09820_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__xor2_2 _09821_ (.A(_04650_),
    .B(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__and4_2 _09822_ (.A(PC[10]),
    .B(PC[11]),
    .C(PC[12]),
    .D(_04475_),
    .X(_04655_));
 sky130_fd_sc_hd__and4_2 _09823_ (.A(PC[13]),
    .B(PC[14]),
    .C(PC[15]),
    .D(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__and4_2 _09824_ (.A(PC[16]),
    .B(PC[17]),
    .C(PC[18]),
    .D(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__and4_2 _09825_ (.A(PC[19]),
    .B(PC[20]),
    .C(PC[21]),
    .D(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__and3_2 _09826_ (.A(PC[22]),
    .B(PC[23]),
    .C(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__and4_2 _09827_ (.A(PC[24]),
    .B(PC[25]),
    .C(PC[26]),
    .D(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__a31o_2 _09828_ (.A1(PC[24]),
    .A2(PC[25]),
    .A3(_04659_),
    .B1(PC[26]),
    .X(_04661_));
 sky130_fd_sc_hd__o211ai_2 _09829_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04661_),
    .C1(_04427_),
    .Y(_04662_));
 sky130_fd_sc_hd__o2bb2ai_2 _09830_ (.A1_N(_04367_),
    .A2_N(_04654_),
    .B1(_04660_),
    .B2(_04662_),
    .Y(\rvsingle.dp.PCNext[26] ));
 sky130_fd_sc_hd__and4_2 _09831_ (.A(PC[25]),
    .B(PC[26]),
    .C(PC[27]),
    .D(_04639_),
    .X(_04663_));
 sky130_fd_sc_hd__a31oi_2 _09832_ (.A1(PC[25]),
    .A2(PC[26]),
    .A3(_04639_),
    .B1(PC[27]),
    .Y(_04664_));
 sky130_fd_sc_hd__or2_2 _09833_ (.A(_04663_),
    .B(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__o21bai_2 _09834_ (.A1(_04618_),
    .A2(PC[26]),
    .B1_N(_04650_),
    .Y(_04666_));
 sky130_fd_sc_hd__xnor2_2 _09835_ (.A(_04617_),
    .B(PC[27]),
    .Y(_04667_));
 sky130_fd_sc_hd__a21o_2 _09836_ (.A1(_04651_),
    .A2(_04666_),
    .B1(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__nand3_2 _09837_ (.A(_04651_),
    .B(_04666_),
    .C(_04667_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand3_2 _09838_ (.A(_04366_),
    .B(_04668_),
    .C(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__o21ai_2 _09839_ (.A1(_04398_),
    .A2(_04665_),
    .B1(_04670_),
    .Y(\rvsingle.dp.PCNext[27] ));
 sky130_fd_sc_hd__or2_2 _09840_ (.A(_04617_),
    .B(PC[28]),
    .X(_04671_));
 sky130_fd_sc_hd__nand2_2 _09841_ (.A(_04617_),
    .B(PC[28]),
    .Y(_04672_));
 sky130_fd_sc_hd__nand2_2 _09842_ (.A(_04671_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__o41a_2 _09843_ (.A1(PC[24]),
    .A2(PC[25]),
    .A3(PC[26]),
    .A4(PC[27]),
    .B1(_04617_),
    .X(_04674_));
 sky130_fd_sc_hd__or4_2 _09844_ (.A(_04644_),
    .B(_04653_),
    .C(_04667_),
    .D(_04634_),
    .X(_04675_));
 sky130_fd_sc_hd__a21oi_2 _09845_ (.A1(_04628_),
    .A2(_04631_),
    .B1(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__nor2_2 _09846_ (.A(_04674_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__xnor2_2 _09847_ (.A(_04673_),
    .B(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__xor2_2 _09848_ (.A(PC[28]),
    .B(_04663_),
    .X(_04679_));
 sky130_fd_sc_hd__o211ai_2 _09849_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04679_),
    .C1(_04427_),
    .Y(_04680_));
 sky130_fd_sc_hd__o21ai_2 _09850_ (.A1(_04678_),
    .A2(_04452_),
    .B1(_04680_),
    .Y(\rvsingle.dp.PCNext[28] ));
 sky130_fd_sc_hd__and3_2 _09851_ (.A(PC[27]),
    .B(PC[28]),
    .C(_04660_),
    .X(_04681_));
 sky130_fd_sc_hd__a21oi_2 _09852_ (.A1(PC[28]),
    .A2(_04663_),
    .B1(PC[29]),
    .Y(_04682_));
 sky130_fd_sc_hd__a21o_2 _09853_ (.A1(PC[29]),
    .A2(_04681_),
    .B1(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__o22a_2 _09854_ (.A1(_04618_),
    .A2(PC[28]),
    .B1(_04674_),
    .B2(_04676_),
    .X(_04684_));
 sky130_fd_sc_hd__a21o_2 _09855_ (.A1(_04618_),
    .A2(PC[28]),
    .B1(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__or2_2 _09856_ (.A(_04617_),
    .B(PC[29]),
    .X(_04686_));
 sky130_fd_sc_hd__nand2_2 _09857_ (.A(_04617_),
    .B(PC[29]),
    .Y(_04687_));
 sky130_fd_sc_hd__nand3_2 _09858_ (.A(_04685_),
    .B(_04686_),
    .C(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__a21o_2 _09859_ (.A1(_04686_),
    .A2(_04687_),
    .B1(_04685_),
    .X(_04689_));
 sky130_fd_sc_hd__nand3_2 _09860_ (.A(_04366_),
    .B(_04688_),
    .C(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__o21ai_2 _09861_ (.A1(_04398_),
    .A2(_04683_),
    .B1(_04690_),
    .Y(\rvsingle.dp.PCNext[29] ));
 sky130_fd_sc_hd__a31oi_2 _09862_ (.A1(PC[28]),
    .A2(PC[29]),
    .A3(_04663_),
    .B1(PC[30]),
    .Y(_04691_));
 sky130_fd_sc_hd__a31o_2 _09863_ (.A1(PC[29]),
    .A2(PC[30]),
    .A3(_04681_),
    .B1(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__nand2_2 _09864_ (.A(_01483_),
    .B(PC[30]),
    .Y(_04693_));
 sky130_fd_sc_hd__or2_2 _09865_ (.A(PC[30]),
    .B(_01483_),
    .X(_04694_));
 sky130_fd_sc_hd__nand4_2 _09866_ (.A(_04671_),
    .B(_04672_),
    .C(_04686_),
    .D(_04687_),
    .Y(_04695_));
 sky130_fd_sc_hd__o21bai_2 _09867_ (.A1(_04674_),
    .A2(_04676_),
    .B1_N(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__o21ai_2 _09868_ (.A1(PC[28]),
    .A2(PC[29]),
    .B1(_04618_),
    .Y(_04697_));
 sky130_fd_sc_hd__a22o_2 _09869_ (.A1(_04693_),
    .A2(_04694_),
    .B1(_04696_),
    .B2(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__nand4_2 _09870_ (.A(_04696_),
    .B(_04697_),
    .C(_04693_),
    .D(_04694_),
    .Y(_04699_));
 sky130_fd_sc_hd__nand3_2 _09871_ (.A(_04366_),
    .B(_04698_),
    .C(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__o21ai_2 _09872_ (.A1(_04398_),
    .A2(_04692_),
    .B1(_04700_),
    .Y(\rvsingle.dp.PCNext[30] ));
 sky130_fd_sc_hd__and2_2 _09873_ (.A(_04618_),
    .B(PC[30]),
    .X(_04701_));
 sky130_fd_sc_hd__or2_2 _09874_ (.A(_04618_),
    .B(PC[31]),
    .X(_04702_));
 sky130_fd_sc_hd__nand2_2 _09875_ (.A(_04618_),
    .B(PC[31]),
    .Y(_04703_));
 sky130_fd_sc_hd__nand4b_2 _09876_ (.A_N(_04701_),
    .B(_04698_),
    .C(_04702_),
    .D(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__a22oi_2 _09877_ (.A1(_04693_),
    .A2(_04694_),
    .B1(_04696_),
    .B2(_04697_),
    .Y(_04705_));
 sky130_fd_sc_hd__nor2_2 _09878_ (.A(_04618_),
    .B(PC[31]),
    .Y(_04706_));
 sky130_fd_sc_hd__and2_2 _09879_ (.A(_04618_),
    .B(PC[31]),
    .X(_04707_));
 sky130_fd_sc_hd__o22ai_2 _09880_ (.A1(_04701_),
    .A2(_04705_),
    .B1(_04706_),
    .B2(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__nand2_2 _09881_ (.A(_04704_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__a41o_2 _09882_ (.A1(PC[28]),
    .A2(PC[29]),
    .A3(PC[30]),
    .A4(_04663_),
    .B1(PC[31]),
    .X(_04710_));
 sky130_fd_sc_hd__nand4_2 _09883_ (.A(PC[29]),
    .B(PC[30]),
    .C(PC[31]),
    .D(_04681_),
    .Y(_04711_));
 sky130_fd_sc_hd__o211ai_2 _09884_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04710_),
    .C1(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__o2bb2ai_2 _09885_ (.A1_N(_04367_),
    .A2_N(_04709_),
    .B1(_04712_),
    .B2(_04365_),
    .Y(\rvsingle.dp.PCNext[31] ));
 sky130_fd_sc_hd__buf_1 _09886_ (.A(_01078_),
    .X(_04713_));
 sky130_fd_sc_hd__and4b_2 _09887_ (.A_N(ReadData[0]),
    .B(_01080_),
    .C(_04121_),
    .D(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__buf_1 _09888_ (.A(_04245_),
    .X(_04715_));
 sky130_fd_sc_hd__a221oi_2 _09889_ (.A1(_04713_),
    .A2(_04715_),
    .B1(_04118_),
    .B2(_04119_),
    .C1(_04129_),
    .Y(_04716_));
 sky130_fd_sc_hd__o32ai_2 _09890_ (.A1(_01169_),
    .A2(_01170_),
    .A3(_02259_),
    .B1(_04714_),
    .B2(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__o21ai_2 _09891_ (.A1(PC[0]),
    .A2(_04426_),
    .B1(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__buf_1 _09892_ (.A(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__buf_1 _09893_ (.A(_04713_),
    .X(_04720_));
 sky130_fd_sc_hd__buf_1 _09894_ (.A(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__buf_1 _09895_ (.A(Instr[11]),
    .X(_04722_));
 sky130_fd_sc_hd__buf_1 _09896_ (.A(Instr[10]),
    .X(_04723_));
 sky130_fd_sc_hd__buf_1 _09897_ (.A(Instr[9]),
    .X(_04724_));
 sky130_fd_sc_hd__nor3_2 _09898_ (.A(_04722_),
    .B(_04723_),
    .C(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__buf_1 _09899_ (.A(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__and2b_2 _09900_ (.A_N(Instr[7]),
    .B(Instr[8]),
    .X(_04727_));
 sky130_fd_sc_hd__buf_1 _09901_ (.A(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__and3_2 _09902_ (.A(_04721_),
    .B(_04726_),
    .C(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__nor2_2 _09903_ (.A(net35),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__a21oi_2 _09904_ (.A1(_04719_),
    .A2(_04729_),
    .B1(_04730_),
    .Y(_00847_));
 sky130_fd_sc_hd__a31o_2 _09905_ (.A1(_04121_),
    .A2(_04713_),
    .A3(ReadData[1]),
    .B1(_04364_),
    .X(_04731_));
 sky130_fd_sc_hd__buf_1 _09906_ (.A(_01069_),
    .X(_04732_));
 sky130_fd_sc_hd__buf_1 _09907_ (.A(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__o31a_2 _09908_ (.A1(_04364_),
    .A2(_04141_),
    .A3(_04733_),
    .B1(DataAdr[1]),
    .X(_04734_));
 sky130_fd_sc_hd__o22a_2 _09909_ (.A1(PC[1]),
    .A2(_04425_),
    .B1(_04731_),
    .B2(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__buf_1 _09910_ (.A(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__buf_1 _09911_ (.A(Instr[7]),
    .X(_04737_));
 sky130_fd_sc_hd__buf_1 _09912_ (.A(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__buf_1 _09913_ (.A(Instr[8]),
    .X(_04739_));
 sky130_fd_sc_hd__or4bb_2 _09914_ (.A(_04738_),
    .B(_04733_),
    .C_N(_04725_),
    .D_N(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__buf_1 _09915_ (.A(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__mux2_2 _09916_ (.A0(_04736_),
    .A1(net798),
    .S(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__buf_1 _09917_ (.A(_04742_),
    .X(_00848_));
 sky130_fd_sc_hd__buf_1 _09918_ (.A(_04140_),
    .X(_04743_));
 sky130_fd_sc_hd__a31o_2 _09919_ (.A1(_04121_),
    .A2(_04713_),
    .A3(ReadData[2]),
    .B1(_04364_),
    .X(_04744_));
 sky130_fd_sc_hd__o31a_2 _09920_ (.A1(_04364_),
    .A2(_04141_),
    .A3(_04732_),
    .B1(DataAdr[2]),
    .X(_04745_));
 sky130_fd_sc_hd__o2bb2a_2 _09921_ (.A1_N(_04397_),
    .A2_N(_04743_),
    .B1(_04744_),
    .B2(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__buf_1 _09922_ (.A(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__mux2_2 _09923_ (.A0(_04747_),
    .A1(\rvsingle.dp.rf.rf[2][2] ),
    .S(_04741_),
    .X(_04748_));
 sky130_fd_sc_hd__buf_1 _09924_ (.A(_04748_),
    .X(_00849_));
 sky130_fd_sc_hd__and3_2 _09925_ (.A(_01080_),
    .B(_04121_),
    .C(_01078_),
    .X(_04749_));
 sky130_fd_sc_hd__buf_1 _09926_ (.A(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__buf_1 _09927_ (.A(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__mux2_2 _09928_ (.A0(DataAdr[3]),
    .A1(ReadData[3]),
    .S(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__nand2_2 _09929_ (.A(_04425_),
    .B(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__o21ai_2 _09930_ (.A1(_04426_),
    .A2(_04406_),
    .B1(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__buf_1 _09931_ (.A(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__mux2_2 _09932_ (.A0(_04755_),
    .A1(\rvsingle.dp.rf.rf[2][3] ),
    .S(_04741_),
    .X(_04756_));
 sky130_fd_sc_hd__buf_1 _09933_ (.A(_04756_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_2 _09934_ (.A0(DataAdr[4]),
    .A1(ReadData[4]),
    .S(_04751_),
    .X(_04757_));
 sky130_fd_sc_hd__and4b_2 _09935_ (.A_N(_04421_),
    .B(_04424_),
    .C(_04505_),
    .D(_04506_),
    .X(_04758_));
 sky130_fd_sc_hd__a21o_2 _09936_ (.A1(_04426_),
    .A2(_04757_),
    .B1(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__buf_1 _09937_ (.A(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__mux2_2 _09938_ (.A0(_04760_),
    .A1(\rvsingle.dp.rf.rf[2][4] ),
    .S(_04741_),
    .X(_04761_));
 sky130_fd_sc_hd__buf_1 _09939_ (.A(_04761_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_2 _09940_ (.A0(DataAdr[5]),
    .A1(ReadData[5]),
    .S(_04751_),
    .X(_04762_));
 sky130_fd_sc_hd__and3_2 _09941_ (.A(_04364_),
    .B(_04430_),
    .C(_04431_),
    .X(_04763_));
 sky130_fd_sc_hd__a21o_2 _09942_ (.A1(_04426_),
    .A2(_04762_),
    .B1(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__buf_1 _09943_ (.A(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__mux2_2 _09944_ (.A0(_04765_),
    .A1(\rvsingle.dp.rf.rf[2][5] ),
    .S(_04741_),
    .X(_04766_));
 sky130_fd_sc_hd__buf_1 _09945_ (.A(_04766_),
    .X(_00852_));
 sky130_fd_sc_hd__or4b_2 _09946_ (.A(_01169_),
    .B(_02259_),
    .C(_01170_),
    .D_N(_04445_),
    .X(_04767_));
 sky130_fd_sc_hd__mux2_2 _09947_ (.A0(DataAdr[6]),
    .A1(ReadData[6]),
    .S(_04751_),
    .X(_04768_));
 sky130_fd_sc_hd__a2bb2o_2 _09948_ (.A1_N(_04767_),
    .A2_N(_04444_),
    .B1(_04426_),
    .B2(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__buf_1 _09949_ (.A(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__mux2_2 _09950_ (.A0(_04770_),
    .A1(\rvsingle.dp.rf.rf[2][6] ),
    .S(_04741_),
    .X(_04771_));
 sky130_fd_sc_hd__buf_1 _09951_ (.A(_04771_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_2 _09952_ (.A0(DataAdr[7]),
    .A1(ReadData[7]),
    .S(_04750_),
    .X(_04772_));
 sky130_fd_sc_hd__mux2_2 _09953_ (.A0(_04772_),
    .A1(_04458_),
    .S(_04743_),
    .X(_04773_));
 sky130_fd_sc_hd__buf_1 _09954_ (.A(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__mux2_2 _09955_ (.A0(_04774_),
    .A1(net406),
    .S(_04741_),
    .X(_04775_));
 sky130_fd_sc_hd__buf_1 _09956_ (.A(_04775_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_2 _09957_ (.A0(DataAdr[8]),
    .A1(ReadData[8]),
    .S(_04751_),
    .X(_04776_));
 sky130_fd_sc_hd__mux2_2 _09958_ (.A0(_04776_),
    .A1(_04468_),
    .S(_04743_),
    .X(_04777_));
 sky130_fd_sc_hd__buf_1 _09959_ (.A(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__mux2_2 _09960_ (.A0(_04778_),
    .A1(net676),
    .S(_04741_),
    .X(_04779_));
 sky130_fd_sc_hd__buf_1 _09961_ (.A(_04779_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_2 _09962_ (.A0(DataAdr[9]),
    .A1(ReadData[9]),
    .S(_04750_),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_2 _09963_ (.A0(_04780_),
    .A1(_04477_),
    .S(_04743_),
    .X(_04781_));
 sky130_fd_sc_hd__buf_1 _09964_ (.A(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__mux2_2 _09965_ (.A0(_04782_),
    .A1(net538),
    .S(_04741_),
    .X(_04783_));
 sky130_fd_sc_hd__buf_1 _09966_ (.A(_04783_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_2 _09967_ (.A0(DataAdr[10]),
    .A1(ReadData[10]),
    .S(_04750_),
    .X(_04784_));
 sky130_fd_sc_hd__mux2_2 _09968_ (.A0(_04784_),
    .A1(_04479_),
    .S(_04743_),
    .X(_04785_));
 sky130_fd_sc_hd__buf_1 _09969_ (.A(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__mux2_2 _09970_ (.A0(_04786_),
    .A1(net570),
    .S(_04741_),
    .X(_04787_));
 sky130_fd_sc_hd__buf_1 _09971_ (.A(_04787_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_2 _09972_ (.A0(DataAdr[11]),
    .A1(ReadData[11]),
    .S(_04750_),
    .X(_04788_));
 sky130_fd_sc_hd__mux2_2 _09973_ (.A0(_04788_),
    .A1(_04502_),
    .S(_04743_),
    .X(_04789_));
 sky130_fd_sc_hd__buf_1 _09974_ (.A(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__buf_1 _09975_ (.A(_04740_),
    .X(_04791_));
 sky130_fd_sc_hd__mux2_2 _09976_ (.A0(_04790_),
    .A1(net339),
    .S(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__buf_1 _09977_ (.A(_04792_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_2 _09978_ (.A0(DataAdr[12]),
    .A1(ReadData[12]),
    .S(_04750_),
    .X(_04793_));
 sky130_fd_sc_hd__mux2_2 _09979_ (.A0(_04793_),
    .A1(_04513_),
    .S(_04364_),
    .X(_04794_));
 sky130_fd_sc_hd__buf_1 _09980_ (.A(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__buf_1 _09981_ (.A(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__mux2_2 _09982_ (.A0(_04796_),
    .A1(net519),
    .S(_04791_),
    .X(_04797_));
 sky130_fd_sc_hd__buf_1 _09983_ (.A(_04797_),
    .X(_00859_));
 sky130_fd_sc_hd__a21oi_2 _09984_ (.A1(_04713_),
    .A2(_04245_),
    .B1(_04268_),
    .Y(_04798_));
 sky130_fd_sc_hd__a31o_2 _09985_ (.A1(ReadData[13]),
    .A2(_04713_),
    .A3(_04245_),
    .B1(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__mux2_2 _09986_ (.A0(_04799_),
    .A1(_04524_),
    .S(_04364_),
    .X(_04800_));
 sky130_fd_sc_hd__buf_1 _09987_ (.A(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__buf_1 _09988_ (.A(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__mux2_2 _09989_ (.A0(_04802_),
    .A1(net648),
    .S(_04791_),
    .X(_04803_));
 sky130_fd_sc_hd__buf_1 _09990_ (.A(_04803_),
    .X(_00860_));
 sky130_fd_sc_hd__o311a_2 _09991_ (.A1(_02909_),
    .A2(_02799_),
    .A3(_02910_),
    .B1(ReadData[14]),
    .C1(_04715_),
    .X(_04804_));
 sky130_fd_sc_hd__a21oi_2 _09992_ (.A1(_02908_),
    .A2(DataAdr[14]),
    .B1(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__or4b_2 _09993_ (.A(_01169_),
    .B(_02259_),
    .C(_01170_),
    .D_N(_04534_),
    .X(_04806_));
 sky130_fd_sc_hd__o21ai_2 _09994_ (.A1(_04365_),
    .A2(_04805_),
    .B1(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__buf_1 _09995_ (.A(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__mux2_2 _09996_ (.A0(_04808_),
    .A1(net602),
    .S(_04791_),
    .X(_04809_));
 sky130_fd_sc_hd__buf_1 _09997_ (.A(_04809_),
    .X(_00861_));
 sky130_fd_sc_hd__o311a_2 _09998_ (.A1(_02909_),
    .A2(_02799_),
    .A3(_02910_),
    .B1(ReadData[15]),
    .C1(_04715_),
    .X(_04810_));
 sky130_fd_sc_hd__a21oi_2 _09999_ (.A1(_04228_),
    .A2(_04396_),
    .B1(_04751_),
    .Y(_04811_));
 sky130_fd_sc_hd__o32a_2 _10000_ (.A1(_01169_),
    .A2(_02259_),
    .A3(_01170_),
    .B1(_04810_),
    .B2(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__a31o_2 _10001_ (.A1(_04505_),
    .A2(_04506_),
    .A3(_04544_),
    .B1(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__buf_1 _10002_ (.A(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__mux2_2 _10003_ (.A0(_04814_),
    .A1(net227),
    .S(_04791_),
    .X(_04815_));
 sky130_fd_sc_hd__buf_1 _10004_ (.A(_04815_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_2 _10005_ (.A0(DataAdr[16]),
    .A1(ReadData[16]),
    .S(_04750_),
    .X(_04816_));
 sky130_fd_sc_hd__mux2_2 _10006_ (.A0(_04816_),
    .A1(_04556_),
    .S(_04743_),
    .X(_04817_));
 sky130_fd_sc_hd__buf_1 _10007_ (.A(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__mux2_2 _10008_ (.A0(_04818_),
    .A1(net403),
    .S(_04791_),
    .X(_04819_));
 sky130_fd_sc_hd__buf_1 _10009_ (.A(_04819_),
    .X(_00863_));
 sky130_fd_sc_hd__or4b_2 _10010_ (.A(_04140_),
    .B(_04141_),
    .C(_04732_),
    .D_N(ReadData[17]),
    .X(_04820_));
 sky130_fd_sc_hd__o21ai_2 _10011_ (.A1(_04751_),
    .A2(_04256_),
    .B1(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__and3_2 _10012_ (.A(_04564_),
    .B(_04565_),
    .C(_04364_),
    .X(_04822_));
 sky130_fd_sc_hd__a21o_2 _10013_ (.A1(_04426_),
    .A2(_04821_),
    .B1(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__buf_1 _10014_ (.A(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__mux2_2 _10015_ (.A0(_04824_),
    .A1(net687),
    .S(_04791_),
    .X(_04825_));
 sky130_fd_sc_hd__buf_1 _10016_ (.A(_04825_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_2 _10017_ (.A0(DataAdr[18]),
    .A1(ReadData[18]),
    .S(_04750_),
    .X(_04826_));
 sky130_fd_sc_hd__mux2_2 _10018_ (.A0(_04826_),
    .A1(_04575_),
    .S(_04743_),
    .X(_04827_));
 sky130_fd_sc_hd__buf_1 _10019_ (.A(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__mux2_2 _10020_ (.A0(_04828_),
    .A1(net524),
    .S(_04791_),
    .X(_04829_));
 sky130_fd_sc_hd__buf_1 _10021_ (.A(_04829_),
    .X(_00865_));
 sky130_fd_sc_hd__or4b_2 _10022_ (.A(_04140_),
    .B(_04141_),
    .C(_04732_),
    .D_N(ReadData[19]),
    .X(_04830_));
 sky130_fd_sc_hd__o21ai_2 _10023_ (.A1(_04751_),
    .A2(_04284_),
    .B1(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__nor2_2 _10024_ (.A(_04425_),
    .B(_04583_),
    .Y(_04832_));
 sky130_fd_sc_hd__a21o_2 _10025_ (.A1(_04425_),
    .A2(_04831_),
    .B1(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__buf_1 _10026_ (.A(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__mux2_2 _10027_ (.A0(_04834_),
    .A1(net615),
    .S(_04791_),
    .X(_04835_));
 sky130_fd_sc_hd__buf_1 _10028_ (.A(_04835_),
    .X(_00866_));
 sky130_fd_sc_hd__o311a_2 _10029_ (.A1(_02909_),
    .A2(_02799_),
    .A3(_02910_),
    .B1(ReadData[20]),
    .C1(_04715_),
    .X(_04836_));
 sky130_fd_sc_hd__a21oi_2 _10030_ (.A1(_02908_),
    .A2(DataAdr[20]),
    .B1(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__and3_2 _10031_ (.A(_04505_),
    .B(_04506_),
    .C(_04595_),
    .X(_04838_));
 sky130_fd_sc_hd__o21bai_2 _10032_ (.A1(_04365_),
    .A2(_04837_),
    .B1_N(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__buf_1 _10033_ (.A(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__mux2_2 _10034_ (.A0(_04840_),
    .A1(net437),
    .S(_04791_),
    .X(_04841_));
 sky130_fd_sc_hd__buf_1 _10035_ (.A(_04841_),
    .X(_00867_));
 sky130_fd_sc_hd__o311a_2 _10036_ (.A1(_02909_),
    .A2(_02799_),
    .A3(_02910_),
    .B1(ReadData[21]),
    .C1(_04715_),
    .X(_04842_));
 sky130_fd_sc_hd__a21oi_2 _10037_ (.A1(_02908_),
    .A2(DataAdr[21]),
    .B1(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__or4_2 _10038_ (.A(_01169_),
    .B(_02259_),
    .C(_01170_),
    .D(_04599_),
    .X(_04844_));
 sky130_fd_sc_hd__o21ai_2 _10039_ (.A1(_04365_),
    .A2(_04843_),
    .B1(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__buf_1 _10040_ (.A(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__buf_1 _10041_ (.A(_04740_),
    .X(_04847_));
 sky130_fd_sc_hd__mux2_2 _10042_ (.A0(_04846_),
    .A1(net605),
    .S(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__buf_1 _10043_ (.A(_04848_),
    .X(_00868_));
 sky130_fd_sc_hd__o311a_2 _10044_ (.A1(_02909_),
    .A2(_02799_),
    .A3(_02910_),
    .B1(ReadData[22]),
    .C1(_04245_),
    .X(_04849_));
 sky130_fd_sc_hd__o21ba_2 _10045_ (.A1(_04751_),
    .A2(_04210_),
    .B1_N(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__or3_2 _10046_ (.A(_01080_),
    .B(_04612_),
    .C(_04613_),
    .X(_04851_));
 sky130_fd_sc_hd__o21ai_2 _10047_ (.A1(_04365_),
    .A2(_04850_),
    .B1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__buf_1 _10048_ (.A(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__mux2_2 _10049_ (.A0(_04853_),
    .A1(net304),
    .S(_04847_),
    .X(_04854_));
 sky130_fd_sc_hd__buf_1 _10050_ (.A(_04854_),
    .X(_00869_));
 sky130_fd_sc_hd__or4b_2 _10051_ (.A(_04140_),
    .B(_04141_),
    .C(_04732_),
    .D_N(ReadData[23]),
    .X(_04855_));
 sky130_fd_sc_hd__nand2_2 _10052_ (.A(_02908_),
    .B(DataAdr[23]),
    .Y(_04856_));
 sky130_fd_sc_hd__a32o_2 _10053_ (.A1(_04505_),
    .A2(_01071_),
    .A3(_01079_),
    .B1(_04855_),
    .B2(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__o21ai_2 _10054_ (.A1(_04426_),
    .A2(_04616_),
    .B1(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__buf_1 _10055_ (.A(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__mux2_2 _10056_ (.A0(_04859_),
    .A1(net582),
    .S(_04847_),
    .X(_04860_));
 sky130_fd_sc_hd__buf_1 _10057_ (.A(_04860_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_2 _10058_ (.A0(DataAdr[24]),
    .A1(ReadData[24]),
    .S(_04750_),
    .X(_04861_));
 sky130_fd_sc_hd__mux2_2 _10059_ (.A0(_04861_),
    .A1(_04641_),
    .S(_04743_),
    .X(_04862_));
 sky130_fd_sc_hd__buf_1 _10060_ (.A(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__mux2_2 _10061_ (.A0(_04863_),
    .A1(net420),
    .S(_04847_),
    .X(_04864_));
 sky130_fd_sc_hd__buf_1 _10062_ (.A(_04864_),
    .X(_00871_));
 sky130_fd_sc_hd__o311a_2 _10063_ (.A1(_02909_),
    .A2(_02799_),
    .A3(_02910_),
    .B1(ReadData[25]),
    .C1(_04245_),
    .X(_04865_));
 sky130_fd_sc_hd__a21o_2 _10064_ (.A1(_02908_),
    .A2(DataAdr[25]),
    .B1(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__nor2_2 _10065_ (.A(_04425_),
    .B(_04643_),
    .Y(_04867_));
 sky130_fd_sc_hd__a21o_2 _10066_ (.A1(_04425_),
    .A2(_04866_),
    .B1(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__buf_1 _10067_ (.A(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__buf_1 _10068_ (.A(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__mux2_2 _10069_ (.A0(_04870_),
    .A1(net759),
    .S(_04847_),
    .X(_04871_));
 sky130_fd_sc_hd__buf_1 _10070_ (.A(_04871_),
    .X(_00872_));
 sky130_fd_sc_hd__o311a_2 _10071_ (.A1(_02909_),
    .A2(_02799_),
    .A3(_02910_),
    .B1(ReadData[26]),
    .C1(_04245_),
    .X(_04872_));
 sky130_fd_sc_hd__a21oi_2 _10072_ (.A1(_02908_),
    .A2(DataAdr[26]),
    .B1(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__or3b_2 _10073_ (.A(_04660_),
    .B(_01080_),
    .C_N(_04661_),
    .X(_04874_));
 sky130_fd_sc_hd__o21ai_2 _10074_ (.A1(_04364_),
    .A2(_04873_),
    .B1(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__buf_1 _10075_ (.A(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__buf_1 _10076_ (.A(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__mux2_2 _10077_ (.A0(_04877_),
    .A1(net223),
    .S(_04847_),
    .X(_04878_));
 sky130_fd_sc_hd__buf_1 _10078_ (.A(_04878_),
    .X(_00873_));
 sky130_fd_sc_hd__buf_1 _10079_ (.A(_02909_),
    .X(_04879_));
 sky130_fd_sc_hd__buf_1 _10080_ (.A(_02799_),
    .X(_04880_));
 sky130_fd_sc_hd__buf_1 _10081_ (.A(_02910_),
    .X(_04881_));
 sky130_fd_sc_hd__o311a_2 _10082_ (.A1(_04879_),
    .A2(_04880_),
    .A3(_04881_),
    .B1(ReadData[27]),
    .C1(_04715_),
    .X(_04882_));
 sky130_fd_sc_hd__a21oi_2 _10083_ (.A1(_02908_),
    .A2(DataAdr[27]),
    .B1(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__nor2_2 _10084_ (.A(_04425_),
    .B(_04665_),
    .Y(_04884_));
 sky130_fd_sc_hd__o21bai_2 _10085_ (.A1(_04365_),
    .A2(_04883_),
    .B1_N(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__buf_1 _10086_ (.A(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__mux2_2 _10087_ (.A0(_04886_),
    .A1(net391),
    .S(_04847_),
    .X(_04887_));
 sky130_fd_sc_hd__buf_1 _10088_ (.A(_04887_),
    .X(_00874_));
 sky130_fd_sc_hd__o311a_2 _10089_ (.A1(_04879_),
    .A2(_04880_),
    .A3(_04881_),
    .B1(ReadData[28]),
    .C1(_04715_),
    .X(_04888_));
 sky130_fd_sc_hd__a21oi_2 _10090_ (.A1(_02908_),
    .A2(DataAdr[28]),
    .B1(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__nand2_2 _10091_ (.A(_04365_),
    .B(_04679_),
    .Y(_04890_));
 sky130_fd_sc_hd__o21ai_2 _10092_ (.A1(_04365_),
    .A2(_04889_),
    .B1(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__buf_1 _10093_ (.A(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__mux2_2 _10094_ (.A0(_04892_),
    .A1(net228),
    .S(_04847_),
    .X(_04893_));
 sky130_fd_sc_hd__buf_1 _10095_ (.A(_04893_),
    .X(_00875_));
 sky130_fd_sc_hd__or4b_2 _10096_ (.A(_04140_),
    .B(_04141_),
    .C(_04732_),
    .D_N(ReadData[29]),
    .X(_04894_));
 sky130_fd_sc_hd__o21ai_2 _10097_ (.A1(_04751_),
    .A2(_04184_),
    .B1(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__nand2_2 _10098_ (.A(_04425_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__o21ai_2 _10099_ (.A1(_04426_),
    .A2(_04683_),
    .B1(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__buf_1 _10100_ (.A(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__mux2_2 _10101_ (.A0(_04898_),
    .A1(net376),
    .S(_04847_),
    .X(_04899_));
 sky130_fd_sc_hd__buf_1 _10102_ (.A(_04899_),
    .X(_00876_));
 sky130_fd_sc_hd__o311a_2 _10103_ (.A1(_04879_),
    .A2(_04880_),
    .A3(_04881_),
    .B1(ReadData[30]),
    .C1(_04715_),
    .X(_04900_));
 sky130_fd_sc_hd__a21oi_2 _10104_ (.A1(_02908_),
    .A2(DataAdr[30]),
    .B1(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__a311o_2 _10105_ (.A1(PC[29]),
    .A2(PC[30]),
    .A3(_04681_),
    .B1(_04691_),
    .C1(_04425_),
    .X(_04902_));
 sky130_fd_sc_hd__o21ai_2 _10106_ (.A1(_04365_),
    .A2(_04901_),
    .B1(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__buf_1 _10107_ (.A(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__mux2_2 _10108_ (.A0(_04904_),
    .A1(net233),
    .S(_04847_),
    .X(_04905_));
 sky130_fd_sc_hd__buf_1 _10109_ (.A(_04905_),
    .X(_00877_));
 sky130_fd_sc_hd__inv_2 _10110_ (.A(net99),
    .Y(_04906_));
 sky130_fd_sc_hd__and3_2 _10111_ (.A(_04711_),
    .B(_04743_),
    .C(_04710_),
    .X(_04907_));
 sky130_fd_sc_hd__buf_1 _10112_ (.A(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__buf_1 _10113_ (.A(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__o311a_2 _10114_ (.A1(_04879_),
    .A2(_04880_),
    .A3(_04881_),
    .B1(ReadData[31]),
    .C1(_04715_),
    .X(_04910_));
 sky130_fd_sc_hd__a22oi_2 _10115_ (.A1(_04713_),
    .A2(_04715_),
    .B1(_04138_),
    .B2(_04132_),
    .Y(_04911_));
 sky130_fd_sc_hd__o32a_2 _10116_ (.A1(_01169_),
    .A2(_02259_),
    .A3(_01170_),
    .B1(_04910_),
    .B2(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__buf_1 _10117_ (.A(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__o21ai_2 _10118_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_04729_),
    .Y(_04914_));
 sky130_fd_sc_hd__o21ai_2 _10119_ (.A1(_04906_),
    .A2(_04729_),
    .B1(_04914_),
    .Y(_00878_));
 sky130_fd_sc_hd__buf_1 _10120_ (.A(_04722_),
    .X(_04915_));
 sky130_fd_sc_hd__buf_1 _10121_ (.A(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__buf_1 _10122_ (.A(_04723_),
    .X(_04917_));
 sky130_fd_sc_hd__buf_1 _10123_ (.A(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__buf_1 _10124_ (.A(Instr[8]),
    .X(_04919_));
 sky130_fd_sc_hd__nor2_2 _10125_ (.A(_04737_),
    .B(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__o31a_2 _10126_ (.A1(_02909_),
    .A2(_02910_),
    .A3(_02799_),
    .B1(_04724_),
    .X(_04921_));
 sky130_fd_sc_hd__buf_1 _10127_ (.A(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__and4_2 _10128_ (.A(_04916_),
    .B(_04918_),
    .C(_04920_),
    .D(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__buf_1 _10129_ (.A(_04920_),
    .X(_04924_));
 sky130_fd_sc_hd__and3_2 _10130_ (.A(_04722_),
    .B(_04723_),
    .C(_04921_),
    .X(_04925_));
 sky130_fd_sc_hd__a21oi_2 _10131_ (.A1(_04924_),
    .A2(_04925_),
    .B1(net24),
    .Y(_04926_));
 sky130_fd_sc_hd__a21oi_2 _10132_ (.A1(_04719_),
    .A2(_04923_),
    .B1(_04926_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_2 _10133_ (.A(_04722_),
    .B(_04723_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand2_2 _10134_ (.A(_04713_),
    .B(_04724_),
    .Y(_04928_));
 sky130_fd_sc_hd__or4_2 _10135_ (.A(_04738_),
    .B(_04739_),
    .C(_04927_),
    .D(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__buf_1 _10136_ (.A(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__mux2_2 _10137_ (.A0(_04736_),
    .A1(\rvsingle.dp.rf.rf[28][1] ),
    .S(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__buf_1 _10138_ (.A(_04931_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_2 _10139_ (.A0(_04747_),
    .A1(net393),
    .S(_04930_),
    .X(_04932_));
 sky130_fd_sc_hd__buf_1 _10140_ (.A(_04932_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_2 _10141_ (.A0(_04755_),
    .A1(\rvsingle.dp.rf.rf[28][3] ),
    .S(_04930_),
    .X(_04933_));
 sky130_fd_sc_hd__buf_1 _10142_ (.A(_04933_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_2 _10143_ (.A0(_04760_),
    .A1(net774),
    .S(_04930_),
    .X(_04934_));
 sky130_fd_sc_hd__buf_1 _10144_ (.A(_04934_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_2 _10145_ (.A0(_04765_),
    .A1(\rvsingle.dp.rf.rf[28][5] ),
    .S(_04930_),
    .X(_04935_));
 sky130_fd_sc_hd__buf_1 _10146_ (.A(_04935_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_2 _10147_ (.A0(_04770_),
    .A1(net656),
    .S(_04930_),
    .X(_04936_));
 sky130_fd_sc_hd__buf_1 _10148_ (.A(_04936_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_2 _10149_ (.A0(_04774_),
    .A1(net809),
    .S(_04930_),
    .X(_04937_));
 sky130_fd_sc_hd__buf_1 _10150_ (.A(_04937_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_2 _10151_ (.A0(_04778_),
    .A1(\rvsingle.dp.rf.rf[28][8] ),
    .S(_04930_),
    .X(_04938_));
 sky130_fd_sc_hd__buf_1 _10152_ (.A(_04938_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_2 _10153_ (.A0(_04782_),
    .A1(net600),
    .S(_04930_),
    .X(_04939_));
 sky130_fd_sc_hd__buf_1 _10154_ (.A(_04939_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_2 _10155_ (.A0(_04786_),
    .A1(\rvsingle.dp.rf.rf[28][10] ),
    .S(_04930_),
    .X(_04940_));
 sky130_fd_sc_hd__buf_1 _10156_ (.A(_04940_),
    .X(_00889_));
 sky130_fd_sc_hd__buf_1 _10157_ (.A(_04929_),
    .X(_04941_));
 sky130_fd_sc_hd__mux2_2 _10158_ (.A0(_04790_),
    .A1(net434),
    .S(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__buf_1 _10159_ (.A(_04942_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_2 _10160_ (.A0(_04796_),
    .A1(net612),
    .S(_04941_),
    .X(_04943_));
 sky130_fd_sc_hd__buf_1 _10161_ (.A(_04943_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_2 _10162_ (.A0(_04802_),
    .A1(net504),
    .S(_04941_),
    .X(_04944_));
 sky130_fd_sc_hd__buf_1 _10163_ (.A(_04944_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_2 _10164_ (.A0(_04808_),
    .A1(net415),
    .S(_04941_),
    .X(_04945_));
 sky130_fd_sc_hd__buf_1 _10165_ (.A(_04945_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_2 _10166_ (.A0(_04814_),
    .A1(\rvsingle.dp.rf.rf[28][15] ),
    .S(_04941_),
    .X(_04946_));
 sky130_fd_sc_hd__buf_1 _10167_ (.A(_04946_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_2 _10168_ (.A0(_04818_),
    .A1(\rvsingle.dp.rf.rf[28][16] ),
    .S(_04941_),
    .X(_04947_));
 sky130_fd_sc_hd__buf_1 _10169_ (.A(_04947_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_2 _10170_ (.A0(_04824_),
    .A1(net755),
    .S(_04941_),
    .X(_04948_));
 sky130_fd_sc_hd__buf_1 _10171_ (.A(_04948_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_2 _10172_ (.A0(_04828_),
    .A1(net707),
    .S(_04941_),
    .X(_04949_));
 sky130_fd_sc_hd__buf_1 _10173_ (.A(_04949_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_2 _10174_ (.A0(_04834_),
    .A1(net732),
    .S(_04941_),
    .X(_04950_));
 sky130_fd_sc_hd__buf_1 _10175_ (.A(_04950_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_2 _10176_ (.A0(_04840_),
    .A1(net273),
    .S(_04941_),
    .X(_04951_));
 sky130_fd_sc_hd__buf_1 _10177_ (.A(_04951_),
    .X(_00899_));
 sky130_fd_sc_hd__buf_1 _10178_ (.A(_04929_),
    .X(_04952_));
 sky130_fd_sc_hd__mux2_2 _10179_ (.A0(_04846_),
    .A1(net279),
    .S(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__buf_1 _10180_ (.A(_04953_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_2 _10181_ (.A0(_04853_),
    .A1(net464),
    .S(_04952_),
    .X(_04954_));
 sky130_fd_sc_hd__buf_1 _10182_ (.A(_04954_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_2 _10183_ (.A0(_04859_),
    .A1(net515),
    .S(_04952_),
    .X(_04955_));
 sky130_fd_sc_hd__buf_1 _10184_ (.A(_04955_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_2 _10185_ (.A0(_04863_),
    .A1(net742),
    .S(_04952_),
    .X(_04956_));
 sky130_fd_sc_hd__buf_1 _10186_ (.A(_04956_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_2 _10187_ (.A0(_04870_),
    .A1(net748),
    .S(_04952_),
    .X(_04957_));
 sky130_fd_sc_hd__buf_1 _10188_ (.A(_04957_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_2 _10189_ (.A0(_04877_),
    .A1(net421),
    .S(_04952_),
    .X(_04958_));
 sky130_fd_sc_hd__buf_1 _10190_ (.A(_04958_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_2 _10191_ (.A0(_04886_),
    .A1(net394),
    .S(_04952_),
    .X(_04959_));
 sky130_fd_sc_hd__buf_1 _10192_ (.A(_04959_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_2 _10193_ (.A0(_04892_),
    .A1(net286),
    .S(_04952_),
    .X(_04960_));
 sky130_fd_sc_hd__buf_1 _10194_ (.A(_04960_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_2 _10195_ (.A0(_04898_),
    .A1(net306),
    .S(_04952_),
    .X(_04961_));
 sky130_fd_sc_hd__buf_1 _10196_ (.A(_04961_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_2 _10197_ (.A0(_04904_),
    .A1(net301),
    .S(_04952_),
    .X(_04962_));
 sky130_fd_sc_hd__buf_1 _10198_ (.A(_04962_),
    .X(_00909_));
 sky130_fd_sc_hd__inv_2 _10199_ (.A(net41),
    .Y(_04963_));
 sky130_fd_sc_hd__o21ai_2 _10200_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_04923_),
    .Y(_04964_));
 sky130_fd_sc_hd__o21ai_2 _10201_ (.A1(_04963_),
    .A2(_04923_),
    .B1(_04964_),
    .Y(_00910_));
 sky130_fd_sc_hd__buf_1 _10202_ (.A(_04724_),
    .X(_04965_));
 sky130_fd_sc_hd__nor2_2 _10203_ (.A(_04965_),
    .B(_04927_),
    .Y(_04966_));
 sky130_fd_sc_hd__buf_1 _10204_ (.A(_04738_),
    .X(_04967_));
 sky130_fd_sc_hd__buf_1 _10205_ (.A(_04739_),
    .X(_04968_));
 sky130_fd_sc_hd__and4_2 _10206_ (.A(_04720_),
    .B(_04966_),
    .C(_04967_),
    .D(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__buf_1 _10207_ (.A(_04966_),
    .X(_04970_));
 sky130_fd_sc_hd__and3_2 _10208_ (.A(_04713_),
    .B(_04919_),
    .C(_04737_),
    .X(_04971_));
 sky130_fd_sc_hd__buf_1 _10209_ (.A(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__buf_1 _10210_ (.A(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__a21oi_2 _10211_ (.A1(_04970_),
    .A2(_04973_),
    .B1(net7),
    .Y(_04974_));
 sky130_fd_sc_hd__a21oi_2 _10212_ (.A1(_04719_),
    .A2(_04969_),
    .B1(_04974_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_2 _10213_ (.A(Instr[7]),
    .B(Instr[8]),
    .Y(_04975_));
 sky130_fd_sc_hd__buf_1 _10214_ (.A(_04732_),
    .X(_04976_));
 sky130_fd_sc_hd__or4_2 _10215_ (.A(_04724_),
    .B(_04927_),
    .C(_04975_),
    .D(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__buf_1 _10216_ (.A(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__mux2_2 _10217_ (.A0(_04736_),
    .A1(net350),
    .S(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__buf_1 _10218_ (.A(_04979_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_2 _10219_ (.A0(_04747_),
    .A1(net639),
    .S(_04978_),
    .X(_04980_));
 sky130_fd_sc_hd__buf_1 _10220_ (.A(_04980_),
    .X(_00913_));
 sky130_fd_sc_hd__buf_1 _10221_ (.A(_04965_),
    .X(_04981_));
 sky130_fd_sc_hd__buf_1 _10222_ (.A(_04915_),
    .X(_04982_));
 sky130_fd_sc_hd__buf_1 _10223_ (.A(_04917_),
    .X(_04983_));
 sky130_fd_sc_hd__and4b_2 _10224_ (.A_N(_04981_),
    .B(_04754_),
    .C(_04982_),
    .D(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__buf_1 _10225_ (.A(_04972_),
    .X(_04985_));
 sky130_fd_sc_hd__a22o_2 _10226_ (.A1(net42),
    .A2(_04978_),
    .B1(_04984_),
    .B2(_04985_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_2 _10227_ (.A0(_04760_),
    .A1(\rvsingle.dp.rf.rf[27][4] ),
    .S(_04978_),
    .X(_04986_));
 sky130_fd_sc_hd__buf_1 _10228_ (.A(_04986_),
    .X(_00915_));
 sky130_fd_sc_hd__and4b_2 _10229_ (.A_N(_04981_),
    .B(_04764_),
    .C(_04982_),
    .D(_04983_),
    .X(_04987_));
 sky130_fd_sc_hd__a22o_2 _10230_ (.A1(net30),
    .A2(_04978_),
    .B1(_04987_),
    .B2(_04985_),
    .X(_00916_));
 sky130_fd_sc_hd__and4b_2 _10231_ (.A_N(_04981_),
    .B(_04769_),
    .C(_04982_),
    .D(_04983_),
    .X(_04988_));
 sky130_fd_sc_hd__a22o_2 _10232_ (.A1(net106),
    .A2(_04978_),
    .B1(_04988_),
    .B2(_04985_),
    .X(_00917_));
 sky130_fd_sc_hd__buf_1 _10233_ (.A(_04977_),
    .X(_04989_));
 sky130_fd_sc_hd__mux2_2 _10234_ (.A0(_04774_),
    .A1(\rvsingle.dp.rf.rf[27][7] ),
    .S(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__buf_1 _10235_ (.A(_04990_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_2 _10236_ (.A0(_04778_),
    .A1(net797),
    .S(_04989_),
    .X(_04991_));
 sky130_fd_sc_hd__buf_1 _10237_ (.A(_04991_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_2 _10238_ (.A0(_04782_),
    .A1(\rvsingle.dp.rf.rf[27][9] ),
    .S(_04989_),
    .X(_04992_));
 sky130_fd_sc_hd__buf_1 _10239_ (.A(_04992_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_2 _10240_ (.A0(_04786_),
    .A1(\rvsingle.dp.rf.rf[27][10] ),
    .S(_04989_),
    .X(_04993_));
 sky130_fd_sc_hd__buf_1 _10241_ (.A(_04993_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_2 _10242_ (.A0(_04790_),
    .A1(\rvsingle.dp.rf.rf[27][11] ),
    .S(_04989_),
    .X(_04994_));
 sky130_fd_sc_hd__buf_1 _10243_ (.A(_04994_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_2 _10244_ (.A0(_04796_),
    .A1(\rvsingle.dp.rf.rf[27][12] ),
    .S(_04989_),
    .X(_04995_));
 sky130_fd_sc_hd__buf_1 _10245_ (.A(_04995_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_2 _10246_ (.A0(_04802_),
    .A1(net763),
    .S(_04989_),
    .X(_04996_));
 sky130_fd_sc_hd__buf_1 _10247_ (.A(_04996_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_2 _10248_ (.A0(_04808_),
    .A1(\rvsingle.dp.rf.rf[27][14] ),
    .S(_04989_),
    .X(_04997_));
 sky130_fd_sc_hd__buf_1 _10249_ (.A(_04997_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_2 _10250_ (.A0(_04814_),
    .A1(net730),
    .S(_04989_),
    .X(_04998_));
 sky130_fd_sc_hd__buf_1 _10251_ (.A(_04998_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_2 _10252_ (.A0(_04818_),
    .A1(net565),
    .S(_04989_),
    .X(_04999_));
 sky130_fd_sc_hd__buf_1 _10253_ (.A(_04999_),
    .X(_00927_));
 sky130_fd_sc_hd__and4b_2 _10254_ (.A_N(_04981_),
    .B(_04823_),
    .C(_04982_),
    .D(_04983_),
    .X(_05000_));
 sky130_fd_sc_hd__a22o_2 _10255_ (.A1(net144),
    .A2(_04978_),
    .B1(_05000_),
    .B2(_04985_),
    .X(_00928_));
 sky130_fd_sc_hd__buf_1 _10256_ (.A(_04977_),
    .X(_05001_));
 sky130_fd_sc_hd__mux2_2 _10257_ (.A0(_04828_),
    .A1(\rvsingle.dp.rf.rf[27][18] ),
    .S(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__buf_1 _10258_ (.A(_05002_),
    .X(_00929_));
 sky130_fd_sc_hd__a31o_2 _10259_ (.A1(_04505_),
    .A2(_01071_),
    .A3(_01062_),
    .B1(_04975_),
    .X(_05003_));
 sky130_fd_sc_hd__buf_1 _10260_ (.A(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__nand2_2 _10261_ (.A(_04834_),
    .B(_04970_),
    .Y(_05005_));
 sky130_fd_sc_hd__a2bb2o_2 _10262_ (.A1_N(_05004_),
    .A2_N(_05005_),
    .B1(_04978_),
    .B2(net156),
    .X(_00930_));
 sky130_fd_sc_hd__and4b_2 _10263_ (.A_N(_04981_),
    .B(_04839_),
    .C(_04982_),
    .D(_04983_),
    .X(_05006_));
 sky130_fd_sc_hd__a22o_2 _10264_ (.A1(net26),
    .A2(_04978_),
    .B1(_05006_),
    .B2(_04985_),
    .X(_00931_));
 sky130_fd_sc_hd__nand2_2 _10265_ (.A(_04846_),
    .B(_04970_),
    .Y(_05007_));
 sky130_fd_sc_hd__a2bb2o_2 _10266_ (.A1_N(_05004_),
    .A2_N(_05007_),
    .B1(_04978_),
    .B2(net154),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_2 _10267_ (.A0(_04853_),
    .A1(\rvsingle.dp.rf.rf[27][22] ),
    .S(_05001_),
    .X(_05008_));
 sky130_fd_sc_hd__buf_1 _10268_ (.A(_05008_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_2 _10269_ (.A0(_04859_),
    .A1(net322),
    .S(_05001_),
    .X(_05009_));
 sky130_fd_sc_hd__buf_1 _10270_ (.A(_05009_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_2 _10271_ (.A0(_04863_),
    .A1(net274),
    .S(_05001_),
    .X(_05010_));
 sky130_fd_sc_hd__buf_1 _10272_ (.A(_05010_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_2 _10273_ (.A0(_04870_),
    .A1(net580),
    .S(_05001_),
    .X(_05011_));
 sky130_fd_sc_hd__buf_1 _10274_ (.A(_05011_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_2 _10275_ (.A0(_04877_),
    .A1(net722),
    .S(_05001_),
    .X(_05012_));
 sky130_fd_sc_hd__buf_1 _10276_ (.A(_05012_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_2 _10277_ (.A0(_04886_),
    .A1(\rvsingle.dp.rf.rf[27][27] ),
    .S(_05001_),
    .X(_05013_));
 sky130_fd_sc_hd__buf_1 _10278_ (.A(_05013_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_2 _10279_ (.A0(_04892_),
    .A1(net289),
    .S(_05001_),
    .X(_05014_));
 sky130_fd_sc_hd__buf_1 _10280_ (.A(_05014_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_2 _10281_ (.A0(_04898_),
    .A1(net710),
    .S(_05001_),
    .X(_05015_));
 sky130_fd_sc_hd__buf_1 _10282_ (.A(_05015_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_2 _10283_ (.A0(_04904_),
    .A1(net272),
    .S(_05001_),
    .X(_05016_));
 sky130_fd_sc_hd__buf_1 _10284_ (.A(_05016_),
    .X(_00941_));
 sky130_fd_sc_hd__inv_2 _10285_ (.A(net68),
    .Y(_05017_));
 sky130_fd_sc_hd__o21ai_2 _10286_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_04969_),
    .Y(_05018_));
 sky130_fd_sc_hd__o21ai_2 _10287_ (.A1(_05017_),
    .A2(_04969_),
    .B1(_05018_),
    .Y(_00942_));
 sky130_fd_sc_hd__and3_2 _10288_ (.A(_04721_),
    .B(_04728_),
    .C(_04966_),
    .X(_05019_));
 sky130_fd_sc_hd__nor2_2 _10289_ (.A(net148),
    .B(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__a21oi_2 _10290_ (.A1(_04719_),
    .A2(_05019_),
    .B1(_05020_),
    .Y(_00943_));
 sky130_fd_sc_hd__or4b_2 _10291_ (.A(_04965_),
    .B(_04927_),
    .C(_04976_),
    .D_N(_04727_),
    .X(_05021_));
 sky130_fd_sc_hd__buf_1 _10292_ (.A(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__mux2_2 _10293_ (.A0(_04736_),
    .A1(net762),
    .S(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__buf_1 _10294_ (.A(_05023_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_2 _10295_ (.A0(_04747_),
    .A1(\rvsingle.dp.rf.rf[26][2] ),
    .S(_05022_),
    .X(_05024_));
 sky130_fd_sc_hd__buf_1 _10296_ (.A(_05024_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_2 _10297_ (.A0(_04755_),
    .A1(net786),
    .S(_05022_),
    .X(_05025_));
 sky130_fd_sc_hd__buf_1 _10298_ (.A(_05025_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_2 _10299_ (.A0(_04760_),
    .A1(net416),
    .S(_05022_),
    .X(_05026_));
 sky130_fd_sc_hd__buf_1 _10300_ (.A(_05026_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_2 _10301_ (.A0(_04765_),
    .A1(net545),
    .S(_05022_),
    .X(_05027_));
 sky130_fd_sc_hd__buf_1 _10302_ (.A(_05027_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_2 _10303_ (.A0(_04770_),
    .A1(net789),
    .S(_05022_),
    .X(_05028_));
 sky130_fd_sc_hd__buf_1 _10304_ (.A(_05028_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_2 _10305_ (.A0(_04774_),
    .A1(\rvsingle.dp.rf.rf[26][7] ),
    .S(_05022_),
    .X(_05029_));
 sky130_fd_sc_hd__buf_1 _10306_ (.A(_05029_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_2 _10307_ (.A0(_04778_),
    .A1(net469),
    .S(_05022_),
    .X(_05030_));
 sky130_fd_sc_hd__buf_1 _10308_ (.A(_05030_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_2 _10309_ (.A0(_04782_),
    .A1(net283),
    .S(_05022_),
    .X(_05031_));
 sky130_fd_sc_hd__buf_1 _10310_ (.A(_05031_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_2 _10311_ (.A0(_04786_),
    .A1(net315),
    .S(_05022_),
    .X(_05032_));
 sky130_fd_sc_hd__buf_1 _10312_ (.A(_05032_),
    .X(_00953_));
 sky130_fd_sc_hd__buf_1 _10313_ (.A(_05021_),
    .X(_05033_));
 sky130_fd_sc_hd__mux2_2 _10314_ (.A0(_04790_),
    .A1(net353),
    .S(_05033_),
    .X(_05034_));
 sky130_fd_sc_hd__buf_1 _10315_ (.A(_05034_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_2 _10316_ (.A0(_04796_),
    .A1(net601),
    .S(_05033_),
    .X(_05035_));
 sky130_fd_sc_hd__buf_1 _10317_ (.A(_05035_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_2 _10318_ (.A0(_04802_),
    .A1(net733),
    .S(_05033_),
    .X(_05036_));
 sky130_fd_sc_hd__buf_1 _10319_ (.A(_05036_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_2 _10320_ (.A0(_04808_),
    .A1(net457),
    .S(_05033_),
    .X(_05037_));
 sky130_fd_sc_hd__buf_1 _10321_ (.A(_05037_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_2 _10322_ (.A0(_04814_),
    .A1(net417),
    .S(_05033_),
    .X(_05038_));
 sky130_fd_sc_hd__buf_1 _10323_ (.A(_05038_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_2 _10324_ (.A0(_04818_),
    .A1(net597),
    .S(_05033_),
    .X(_05039_));
 sky130_fd_sc_hd__buf_1 _10325_ (.A(_05039_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_2 _10326_ (.A0(_04824_),
    .A1(net573),
    .S(_05033_),
    .X(_05040_));
 sky130_fd_sc_hd__buf_1 _10327_ (.A(_05040_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_2 _10328_ (.A0(_04828_),
    .A1(net418),
    .S(_05033_),
    .X(_05041_));
 sky130_fd_sc_hd__buf_1 _10329_ (.A(_05041_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_2 _10330_ (.A0(_04834_),
    .A1(\rvsingle.dp.rf.rf[26][19] ),
    .S(_05033_),
    .X(_05042_));
 sky130_fd_sc_hd__buf_1 _10331_ (.A(_05042_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_2 _10332_ (.A0(_04840_),
    .A1(net718),
    .S(_05033_),
    .X(_05043_));
 sky130_fd_sc_hd__buf_1 _10333_ (.A(_05043_),
    .X(_00963_));
 sky130_fd_sc_hd__buf_1 _10334_ (.A(_05021_),
    .X(_05044_));
 sky130_fd_sc_hd__mux2_2 _10335_ (.A0(_04846_),
    .A1(net366),
    .S(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__buf_1 _10336_ (.A(_05045_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_2 _10337_ (.A0(_04853_),
    .A1(net456),
    .S(_05044_),
    .X(_05046_));
 sky130_fd_sc_hd__buf_1 _10338_ (.A(_05046_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_2 _10339_ (.A0(_04859_),
    .A1(net320),
    .S(_05044_),
    .X(_05047_));
 sky130_fd_sc_hd__buf_1 _10340_ (.A(_05047_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_2 _10341_ (.A0(_04863_),
    .A1(net229),
    .S(_05044_),
    .X(_05048_));
 sky130_fd_sc_hd__buf_1 _10342_ (.A(_05048_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_2 _10343_ (.A0(_04870_),
    .A1(net425),
    .S(_05044_),
    .X(_05049_));
 sky130_fd_sc_hd__buf_1 _10344_ (.A(_05049_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_2 _10345_ (.A0(_04877_),
    .A1(net405),
    .S(_05044_),
    .X(_05050_));
 sky130_fd_sc_hd__buf_1 _10346_ (.A(_05050_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_2 _10347_ (.A0(_04886_),
    .A1(net382),
    .S(_05044_),
    .X(_05051_));
 sky130_fd_sc_hd__buf_1 _10348_ (.A(_05051_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_2 _10349_ (.A0(_04892_),
    .A1(net297),
    .S(_05044_),
    .X(_05052_));
 sky130_fd_sc_hd__buf_1 _10350_ (.A(_05052_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_2 _10351_ (.A0(_04898_),
    .A1(net446),
    .S(_05044_),
    .X(_05053_));
 sky130_fd_sc_hd__buf_1 _10352_ (.A(_05053_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_2 _10353_ (.A0(_04904_),
    .A1(net337),
    .S(_05044_),
    .X(_05054_));
 sky130_fd_sc_hd__buf_1 _10354_ (.A(_05054_),
    .X(_00973_));
 sky130_fd_sc_hd__inv_2 _10355_ (.A(net84),
    .Y(_05055_));
 sky130_fd_sc_hd__o21ai_2 _10356_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_05019_),
    .Y(_05056_));
 sky130_fd_sc_hd__o21ai_2 _10357_ (.A1(_05055_),
    .A2(_05019_),
    .B1(_05056_),
    .Y(_00974_));
 sky130_fd_sc_hd__nor2b_2 _10358_ (.A(_04919_),
    .B_N(Instr[7]),
    .Y(_05057_));
 sky130_fd_sc_hd__buf_1 _10359_ (.A(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__and3_2 _10360_ (.A(_04721_),
    .B(_04970_),
    .C(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__buf_1 _10361_ (.A(_04720_),
    .X(_05060_));
 sky130_fd_sc_hd__buf_1 _10362_ (.A(_05057_),
    .X(_05061_));
 sky130_fd_sc_hd__a31o_2 _10363_ (.A1(_05060_),
    .A2(_04970_),
    .A3(_05061_),
    .B1(net581),
    .X(_05062_));
 sky130_fd_sc_hd__a21boi_2 _10364_ (.A1(_04719_),
    .A2(_05059_),
    .B1_N(_05062_),
    .Y(_00975_));
 sky130_fd_sc_hd__or3b_2 _10365_ (.A(Instr[8]),
    .B(_04732_),
    .C_N(Instr[7]),
    .X(_05063_));
 sky130_fd_sc_hd__or3_2 _10366_ (.A(_04965_),
    .B(_04927_),
    .C(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__buf_1 _10367_ (.A(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__mux2_2 _10368_ (.A0(_04736_),
    .A1(net370),
    .S(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__buf_1 _10369_ (.A(_05066_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_2 _10370_ (.A0(_04747_),
    .A1(net659),
    .S(_05065_),
    .X(_05067_));
 sky130_fd_sc_hd__buf_1 _10371_ (.A(_05067_),
    .X(_00977_));
 sky130_fd_sc_hd__buf_1 _10372_ (.A(_05058_),
    .X(_05068_));
 sky130_fd_sc_hd__buf_1 _10373_ (.A(_05060_),
    .X(_05069_));
 sky130_fd_sc_hd__a32o_2 _10374_ (.A1(_04984_),
    .A2(_05068_),
    .A3(_05069_),
    .B1(_05065_),
    .B2(net5),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_2 _10375_ (.A0(_04760_),
    .A1(net586),
    .S(_05065_),
    .X(_05070_));
 sky130_fd_sc_hd__buf_1 _10376_ (.A(_05070_),
    .X(_00979_));
 sky130_fd_sc_hd__a32o_2 _10377_ (.A1(_04987_),
    .A2(_05068_),
    .A3(_05069_),
    .B1(_05065_),
    .B2(net2),
    .X(_00980_));
 sky130_fd_sc_hd__a32o_2 _10378_ (.A1(_04988_),
    .A2(_05068_),
    .A3(_05069_),
    .B1(_05065_),
    .B2(net75),
    .X(_00981_));
 sky130_fd_sc_hd__buf_1 _10379_ (.A(_05064_),
    .X(_05071_));
 sky130_fd_sc_hd__mux2_2 _10380_ (.A0(_04774_),
    .A1(net389),
    .S(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__buf_1 _10381_ (.A(_05072_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_2 _10382_ (.A0(_04778_),
    .A1(\rvsingle.dp.rf.rf[25][8] ),
    .S(_05071_),
    .X(_05073_));
 sky130_fd_sc_hd__buf_1 _10383_ (.A(_05073_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_2 _10384_ (.A0(_04782_),
    .A1(net787),
    .S(_05071_),
    .X(_05074_));
 sky130_fd_sc_hd__buf_1 _10385_ (.A(_05074_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_2 _10386_ (.A0(_04786_),
    .A1(\rvsingle.dp.rf.rf[25][10] ),
    .S(_05071_),
    .X(_05075_));
 sky130_fd_sc_hd__buf_1 _10387_ (.A(_05075_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_2 _10388_ (.A0(_04790_),
    .A1(\rvsingle.dp.rf.rf[25][11] ),
    .S(_05071_),
    .X(_05076_));
 sky130_fd_sc_hd__buf_1 _10389_ (.A(_05076_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_2 _10390_ (.A0(_04796_),
    .A1(net764),
    .S(_05071_),
    .X(_05077_));
 sky130_fd_sc_hd__buf_1 _10391_ (.A(_05077_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_2 _10392_ (.A0(_04802_),
    .A1(net818),
    .S(_05071_),
    .X(_05078_));
 sky130_fd_sc_hd__buf_1 _10393_ (.A(_05078_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_2 _10394_ (.A0(_04808_),
    .A1(net523),
    .S(_05071_),
    .X(_05079_));
 sky130_fd_sc_hd__buf_1 _10395_ (.A(_05079_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_2 _10396_ (.A0(_04814_),
    .A1(net480),
    .S(_05071_),
    .X(_05080_));
 sky130_fd_sc_hd__buf_1 _10397_ (.A(_05080_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_2 _10398_ (.A0(_04818_),
    .A1(net343),
    .S(_05071_),
    .X(_05081_));
 sky130_fd_sc_hd__buf_1 _10399_ (.A(_05081_),
    .X(_00991_));
 sky130_fd_sc_hd__a32o_2 _10400_ (.A1(_05000_),
    .A2(_05068_),
    .A3(_05069_),
    .B1(_05065_),
    .B2(net10),
    .X(_00992_));
 sky130_fd_sc_hd__buf_1 _10401_ (.A(_05064_),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_2 _10402_ (.A0(_04828_),
    .A1(\rvsingle.dp.rf.rf[25][18] ),
    .S(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__buf_1 _10403_ (.A(_05083_),
    .X(_00993_));
 sky130_fd_sc_hd__buf_1 _10404_ (.A(_05063_),
    .X(_05084_));
 sky130_fd_sc_hd__buf_1 _10405_ (.A(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__a2bb2o_2 _10406_ (.A1_N(_05005_),
    .A2_N(_05085_),
    .B1(_05065_),
    .B2(net146),
    .X(_00994_));
 sky130_fd_sc_hd__a32o_2 _10407_ (.A1(_05006_),
    .A2(_05068_),
    .A3(_05069_),
    .B1(_05065_),
    .B2(net6),
    .X(_00995_));
 sky130_fd_sc_hd__a2bb2o_2 _10408_ (.A1_N(_05007_),
    .A2_N(_05085_),
    .B1(_05065_),
    .B2(net130),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_2 _10409_ (.A0(_04853_),
    .A1(net234),
    .S(_05082_),
    .X(_05086_));
 sky130_fd_sc_hd__buf_1 _10410_ (.A(_05086_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_2 _10411_ (.A0(_04859_),
    .A1(net245),
    .S(_05082_),
    .X(_05087_));
 sky130_fd_sc_hd__buf_1 _10412_ (.A(_05087_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_2 _10413_ (.A0(_04863_),
    .A1(net308),
    .S(_05082_),
    .X(_05088_));
 sky130_fd_sc_hd__buf_1 _10414_ (.A(_05088_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_2 _10415_ (.A0(_04870_),
    .A1(net496),
    .S(_05082_),
    .X(_05089_));
 sky130_fd_sc_hd__buf_1 _10416_ (.A(_05089_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_2 _10417_ (.A0(_04877_),
    .A1(net769),
    .S(_05082_),
    .X(_05090_));
 sky130_fd_sc_hd__buf_1 _10418_ (.A(_05090_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_2 _10419_ (.A0(_04886_),
    .A1(net693),
    .S(_05082_),
    .X(_05091_));
 sky130_fd_sc_hd__buf_1 _10420_ (.A(_05091_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_2 _10421_ (.A0(_04892_),
    .A1(net236),
    .S(_05082_),
    .X(_05092_));
 sky130_fd_sc_hd__buf_1 _10422_ (.A(_05092_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_2 _10423_ (.A0(_04898_),
    .A1(net616),
    .S(_05082_),
    .X(_05093_));
 sky130_fd_sc_hd__buf_1 _10424_ (.A(_05093_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_2 _10425_ (.A0(_04904_),
    .A1(net371),
    .S(_05082_),
    .X(_05094_));
 sky130_fd_sc_hd__buf_1 _10426_ (.A(_05094_),
    .X(_01005_));
 sky130_fd_sc_hd__inv_2 _10427_ (.A(net67),
    .Y(_05095_));
 sky130_fd_sc_hd__o21ai_2 _10428_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_05059_),
    .Y(_05096_));
 sky130_fd_sc_hd__o21ai_2 _10429_ (.A1(_05095_),
    .A2(_05059_),
    .B1(_05096_),
    .Y(_01006_));
 sky130_fd_sc_hd__buf_1 _10430_ (.A(_04720_),
    .X(_05097_));
 sky130_fd_sc_hd__and3_2 _10431_ (.A(_05097_),
    .B(_04924_),
    .C(_04970_),
    .X(_05098_));
 sky130_fd_sc_hd__o31a_2 _10432_ (.A1(_04879_),
    .A2(_04881_),
    .A3(_04880_),
    .B1(_04920_),
    .X(_05099_));
 sky130_fd_sc_hd__a21oi_2 _10433_ (.A1(_04970_),
    .A2(_05099_),
    .B1(net17),
    .Y(_05100_));
 sky130_fd_sc_hd__a21oi_2 _10434_ (.A1(_04719_),
    .A2(_05098_),
    .B1(_05100_),
    .Y(_01007_));
 sky130_fd_sc_hd__or2_2 _10435_ (.A(_04724_),
    .B(_04927_),
    .X(_05101_));
 sky130_fd_sc_hd__or4_2 _10436_ (.A(_04737_),
    .B(_04919_),
    .C(_04733_),
    .D(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__buf_1 _10437_ (.A(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__mux2_2 _10438_ (.A0(_04736_),
    .A1(net771),
    .S(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__buf_1 _10439_ (.A(_05104_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_2 _10440_ (.A0(_04747_),
    .A1(\rvsingle.dp.rf.rf[24][2] ),
    .S(_05103_),
    .X(_05105_));
 sky130_fd_sc_hd__buf_1 _10441_ (.A(_05105_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_2 _10442_ (.A0(_04755_),
    .A1(net731),
    .S(_05103_),
    .X(_05106_));
 sky130_fd_sc_hd__buf_1 _10443_ (.A(_05106_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_2 _10444_ (.A0(_04760_),
    .A1(net445),
    .S(_05103_),
    .X(_05107_));
 sky130_fd_sc_hd__buf_1 _10445_ (.A(_05107_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_2 _10446_ (.A0(_04765_),
    .A1(net765),
    .S(_05103_),
    .X(_05108_));
 sky130_fd_sc_hd__buf_1 _10447_ (.A(_05108_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_2 _10448_ (.A0(_04770_),
    .A1(\rvsingle.dp.rf.rf[24][6] ),
    .S(_05103_),
    .X(_05109_));
 sky130_fd_sc_hd__buf_1 _10449_ (.A(_05109_),
    .X(_01013_));
 sky130_fd_sc_hd__buf_1 _10450_ (.A(_05102_),
    .X(_05110_));
 sky130_fd_sc_hd__mux2_2 _10451_ (.A0(_04774_),
    .A1(\rvsingle.dp.rf.rf[24][7] ),
    .S(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__buf_1 _10452_ (.A(_05111_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_2 _10453_ (.A0(_04778_),
    .A1(\rvsingle.dp.rf.rf[24][8] ),
    .S(_05110_),
    .X(_05112_));
 sky130_fd_sc_hd__buf_1 _10454_ (.A(_05112_),
    .X(_01015_));
 sky130_fd_sc_hd__buf_1 _10455_ (.A(_04879_),
    .X(_05113_));
 sky130_fd_sc_hd__buf_1 _10456_ (.A(_04881_),
    .X(_05114_));
 sky130_fd_sc_hd__buf_1 _10457_ (.A(_04880_),
    .X(_05115_));
 sky130_fd_sc_hd__o311a_2 _10458_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_04924_),
    .C1(_04781_),
    .X(_05116_));
 sky130_fd_sc_hd__a22o_2 _10459_ (.A1(net8),
    .A2(_05103_),
    .B1(_05116_),
    .B2(_04970_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_2 _10460_ (.A0(_04786_),
    .A1(\rvsingle.dp.rf.rf[24][10] ),
    .S(_05110_),
    .X(_05117_));
 sky130_fd_sc_hd__buf_1 _10461_ (.A(_05117_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_2 _10462_ (.A0(_04790_),
    .A1(\rvsingle.dp.rf.rf[24][11] ),
    .S(_05110_),
    .X(_05118_));
 sky130_fd_sc_hd__buf_1 _10463_ (.A(_05118_),
    .X(_01018_));
 sky130_fd_sc_hd__o311a_2 _10464_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_04924_),
    .C1(_04795_),
    .X(_05119_));
 sky130_fd_sc_hd__a22o_2 _10465_ (.A1(net166),
    .A2(_05103_),
    .B1(_05119_),
    .B2(_04970_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_2 _10466_ (.A0(_04802_),
    .A1(\rvsingle.dp.rf.rf[24][13] ),
    .S(_05110_),
    .X(_05120_));
 sky130_fd_sc_hd__buf_1 _10467_ (.A(_05120_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_2 _10468_ (.A0(_04808_),
    .A1(\rvsingle.dp.rf.rf[24][14] ),
    .S(_05110_),
    .X(_05121_));
 sky130_fd_sc_hd__buf_1 _10469_ (.A(_05121_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_2 _10470_ (.A0(_04814_),
    .A1(\rvsingle.dp.rf.rf[24][15] ),
    .S(_05110_),
    .X(_05122_));
 sky130_fd_sc_hd__buf_1 _10471_ (.A(_05122_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_2 _10472_ (.A0(_04818_),
    .A1(net237),
    .S(_05110_),
    .X(_05123_));
 sky130_fd_sc_hd__buf_1 _10473_ (.A(_05123_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_2 _10474_ (.A0(_04824_),
    .A1(net738),
    .S(_05110_),
    .X(_05124_));
 sky130_fd_sc_hd__buf_1 _10475_ (.A(_05124_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_2 _10476_ (.A0(_04828_),
    .A1(net539),
    .S(_05110_),
    .X(_05125_));
 sky130_fd_sc_hd__buf_1 _10477_ (.A(_05125_),
    .X(_01025_));
 sky130_fd_sc_hd__buf_1 _10478_ (.A(_05102_),
    .X(_05126_));
 sky130_fd_sc_hd__mux2_2 _10479_ (.A0(_04834_),
    .A1(net625),
    .S(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__buf_1 _10480_ (.A(_05127_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_2 _10481_ (.A0(_04840_),
    .A1(net626),
    .S(_05126_),
    .X(_05128_));
 sky130_fd_sc_hd__buf_1 _10482_ (.A(_05128_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_2 _10483_ (.A0(_04846_),
    .A1(net436),
    .S(_05126_),
    .X(_05129_));
 sky130_fd_sc_hd__buf_1 _10484_ (.A(_05129_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_2 _10485_ (.A0(_04853_),
    .A1(net770),
    .S(_05126_),
    .X(_05130_));
 sky130_fd_sc_hd__buf_1 _10486_ (.A(_05130_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_2 _10487_ (.A0(_04859_),
    .A1(net528),
    .S(_05126_),
    .X(_05131_));
 sky130_fd_sc_hd__buf_1 _10488_ (.A(_05131_),
    .X(_01030_));
 sky130_fd_sc_hd__buf_1 _10489_ (.A(_04862_),
    .X(_05132_));
 sky130_fd_sc_hd__o311a_2 _10490_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_04924_),
    .C1(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__a22o_2 _10491_ (.A1(net23),
    .A2(_05103_),
    .B1(_05133_),
    .B2(_04970_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_2 _10492_ (.A0(_04870_),
    .A1(net678),
    .S(_05126_),
    .X(_05134_));
 sky130_fd_sc_hd__buf_1 _10493_ (.A(_05134_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_2 _10494_ (.A0(_04877_),
    .A1(net462),
    .S(_05126_),
    .X(_05135_));
 sky130_fd_sc_hd__buf_1 _10495_ (.A(_05135_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_2 _10496_ (.A0(_04886_),
    .A1(net453),
    .S(_05126_),
    .X(_05136_));
 sky130_fd_sc_hd__buf_1 _10497_ (.A(_05136_),
    .X(_01034_));
 sky130_fd_sc_hd__nand2_2 _10498_ (.A(_04892_),
    .B(_05099_),
    .Y(_05137_));
 sky130_fd_sc_hd__a2bb2o_2 _10499_ (.A1_N(_05101_),
    .A2_N(_05137_),
    .B1(_05103_),
    .B2(net216),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_2 _10500_ (.A0(_04898_),
    .A1(net341),
    .S(_05126_),
    .X(_05138_));
 sky130_fd_sc_hd__buf_1 _10501_ (.A(_05138_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_2 _10502_ (.A0(_04904_),
    .A1(net323),
    .S(_05126_),
    .X(_05139_));
 sky130_fd_sc_hd__buf_1 _10503_ (.A(_05139_),
    .X(_01037_));
 sky130_fd_sc_hd__inv_2 _10504_ (.A(net77),
    .Y(_05140_));
 sky130_fd_sc_hd__o21ai_2 _10505_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_05098_),
    .Y(_05141_));
 sky130_fd_sc_hd__o21ai_2 _10506_ (.A1(_05140_),
    .A2(_05098_),
    .B1(_05141_),
    .Y(_01038_));
 sky130_fd_sc_hd__nor3b_2 _10507_ (.A(_04915_),
    .B(_04965_),
    .C_N(_04917_),
    .Y(_05142_));
 sky130_fd_sc_hd__and3_2 _10508_ (.A(_05097_),
    .B(_05058_),
    .C(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__o31a_2 _10509_ (.A1(_04879_),
    .A2(_04881_),
    .A3(_04880_),
    .B1(_05057_),
    .X(_05144_));
 sky130_fd_sc_hd__buf_1 _10510_ (.A(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__buf_1 _10511_ (.A(_05142_),
    .X(_05146_));
 sky130_fd_sc_hd__a21oi_2 _10512_ (.A1(_05145_),
    .A2(_05146_),
    .B1(net1),
    .Y(_05147_));
 sky130_fd_sc_hd__a21oi_2 _10513_ (.A1(_04719_),
    .A2(_05143_),
    .B1(_05147_),
    .Y(_01039_));
 sky130_fd_sc_hd__or3b_2 _10514_ (.A(Instr[11]),
    .B(_04724_),
    .C_N(Instr[10]),
    .X(_05148_));
 sky130_fd_sc_hd__buf_1 _10515_ (.A(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__or4b_2 _10516_ (.A(Instr[8]),
    .B(_04732_),
    .C(_05149_),
    .D_N(Instr[7]),
    .X(_05150_));
 sky130_fd_sc_hd__buf_1 _10517_ (.A(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__buf_1 _10518_ (.A(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__mux2_2 _10519_ (.A0(_04736_),
    .A1(\rvsingle.dp.rf.rf[9][1] ),
    .S(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__buf_1 _10520_ (.A(_05153_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_2 _10521_ (.A0(_04747_),
    .A1(\rvsingle.dp.rf.rf[9][2] ),
    .S(_05152_),
    .X(_05154_));
 sky130_fd_sc_hd__buf_1 _10522_ (.A(_05154_),
    .X(_01041_));
 sky130_fd_sc_hd__buf_1 _10523_ (.A(_05152_),
    .X(_05155_));
 sky130_fd_sc_hd__o311a_2 _10524_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_05061_),
    .C1(_04754_),
    .X(_05156_));
 sky130_fd_sc_hd__buf_1 _10525_ (.A(_05146_),
    .X(_05157_));
 sky130_fd_sc_hd__a22o_2 _10526_ (.A1(net150),
    .A2(_05155_),
    .B1(_05156_),
    .B2(_05157_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_2 _10527_ (.A0(_04760_),
    .A1(net671),
    .S(_05152_),
    .X(_05158_));
 sky130_fd_sc_hd__buf_1 _10528_ (.A(_05158_),
    .X(_01043_));
 sky130_fd_sc_hd__o311a_2 _10529_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_05061_),
    .C1(_04764_),
    .X(_05159_));
 sky130_fd_sc_hd__a22o_2 _10530_ (.A1(net88),
    .A2(_05155_),
    .B1(_05159_),
    .B2(_05157_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_2 _10531_ (.A0(_04770_),
    .A1(net768),
    .S(_05152_),
    .X(_05160_));
 sky130_fd_sc_hd__buf_1 _10532_ (.A(_05160_),
    .X(_01045_));
 sky130_fd_sc_hd__o311a_2 _10533_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_05061_),
    .C1(_04773_),
    .X(_05161_));
 sky130_fd_sc_hd__a22o_2 _10534_ (.A1(net78),
    .A2(_05155_),
    .B1(_05161_),
    .B2(_05157_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_2 _10535_ (.A0(_04778_),
    .A1(\rvsingle.dp.rf.rf[9][8] ),
    .S(_05152_),
    .X(_05162_));
 sky130_fd_sc_hd__buf_1 _10536_ (.A(_05162_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_2 _10537_ (.A0(_04782_),
    .A1(net312),
    .S(_05152_),
    .X(_05163_));
 sky130_fd_sc_hd__buf_1 _10538_ (.A(_05163_),
    .X(_01048_));
 sky130_fd_sc_hd__o311a_2 _10539_ (.A1(_04879_),
    .A2(_04881_),
    .A3(_04880_),
    .B1(_05061_),
    .C1(_04785_),
    .X(_05164_));
 sky130_fd_sc_hd__a22o_2 _10540_ (.A1(net50),
    .A2(_05155_),
    .B1(_05164_),
    .B2(_05157_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_2 _10541_ (.A0(_04790_),
    .A1(net767),
    .S(_05152_),
    .X(_05165_));
 sky130_fd_sc_hd__buf_1 _10542_ (.A(_05165_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_2 _10543_ (.A0(_04796_),
    .A1(net592),
    .S(_05151_),
    .X(_05166_));
 sky130_fd_sc_hd__buf_1 _10544_ (.A(_05166_),
    .X(_01051_));
 sky130_fd_sc_hd__buf_1 _10545_ (.A(_05149_),
    .X(_05167_));
 sky130_fd_sc_hd__nand2_2 _10546_ (.A(_04802_),
    .B(_05145_),
    .Y(_05168_));
 sky130_fd_sc_hd__a2bb2o_2 _10547_ (.A1_N(_05167_),
    .A2_N(_05168_),
    .B1(_05155_),
    .B2(net114),
    .X(_01052_));
 sky130_fd_sc_hd__nand2_2 _10548_ (.A(_04808_),
    .B(_05144_),
    .Y(_05169_));
 sky130_fd_sc_hd__a2bb2o_2 _10549_ (.A1_N(_05167_),
    .A2_N(_05169_),
    .B1(_05155_),
    .B2(net139),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_2 _10550_ (.A0(_04814_),
    .A1(net372),
    .S(_05151_),
    .X(_05170_));
 sky130_fd_sc_hd__buf_1 _10551_ (.A(_05170_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_2 _10552_ (.A0(_04818_),
    .A1(net664),
    .S(_05151_),
    .X(_05171_));
 sky130_fd_sc_hd__buf_1 _10553_ (.A(_05171_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_2 _10554_ (.A0(_04824_),
    .A1(net478),
    .S(_05151_),
    .X(_05172_));
 sky130_fd_sc_hd__buf_1 _10555_ (.A(_05172_),
    .X(_01056_));
 sky130_fd_sc_hd__buf_1 _10556_ (.A(_04827_),
    .X(_05173_));
 sky130_fd_sc_hd__o311a_2 _10557_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_05061_),
    .C1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__a22o_2 _10558_ (.A1(net155),
    .A2(_05155_),
    .B1(_05174_),
    .B2(_05157_),
    .X(_01057_));
 sky130_fd_sc_hd__nand2_2 _10559_ (.A(_04834_),
    .B(_05145_),
    .Y(_05175_));
 sky130_fd_sc_hd__a2bb2o_2 _10560_ (.A1_N(_05167_),
    .A2_N(_05175_),
    .B1(_05155_),
    .B2(net94),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_2 _10561_ (.A0(_04840_),
    .A1(net669),
    .S(_05151_),
    .X(_05176_));
 sky130_fd_sc_hd__buf_1 _10562_ (.A(_05176_),
    .X(_00033_));
 sky130_fd_sc_hd__nand2_2 _10563_ (.A(_04846_),
    .B(_05144_),
    .Y(_05177_));
 sky130_fd_sc_hd__a2bb2o_2 _10564_ (.A1_N(_05167_),
    .A2_N(_05177_),
    .B1(_05155_),
    .B2(net186),
    .X(_00034_));
 sky130_fd_sc_hd__o311a_2 _10565_ (.A1(_04879_),
    .A2(_04881_),
    .A3(_04880_),
    .B1(_05058_),
    .C1(_04852_),
    .X(_05178_));
 sky130_fd_sc_hd__a22o_2 _10566_ (.A1(net27),
    .A2(_05155_),
    .B1(_05178_),
    .B2(_05157_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_2 _10567_ (.A0(_04859_),
    .A1(\rvsingle.dp.rf.rf[9][23] ),
    .S(_05151_),
    .X(_05179_));
 sky130_fd_sc_hd__buf_1 _10568_ (.A(_05179_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_2 _10569_ (.A0(_04863_),
    .A1(net254),
    .S(_05151_),
    .X(_05180_));
 sky130_fd_sc_hd__buf_1 _10570_ (.A(_05180_),
    .X(_00037_));
 sky130_fd_sc_hd__o311a_2 _10571_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_05061_),
    .C1(_04869_),
    .X(_05181_));
 sky130_fd_sc_hd__a22o_2 _10572_ (.A1(net66),
    .A2(_05152_),
    .B1(_05181_),
    .B2(_05157_),
    .X(_00038_));
 sky130_fd_sc_hd__o311a_2 _10573_ (.A1(_04879_),
    .A2(_04881_),
    .A3(_04880_),
    .B1(_05058_),
    .C1(_04876_),
    .X(_05182_));
 sky130_fd_sc_hd__a22o_2 _10574_ (.A1(net214),
    .A2(_05152_),
    .B1(_05182_),
    .B2(_05157_),
    .X(_00039_));
 sky130_fd_sc_hd__buf_1 _10575_ (.A(_05144_),
    .X(_05183_));
 sky130_fd_sc_hd__a21oi_2 _10576_ (.A1(_05145_),
    .A2(_05146_),
    .B1(_03924_),
    .Y(_05184_));
 sky130_fd_sc_hd__a31o_2 _10577_ (.A1(_04886_),
    .A2(_05183_),
    .A3(_05146_),
    .B1(_05184_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_2 _10578_ (.A0(_04892_),
    .A1(net294),
    .S(_05151_),
    .X(_05185_));
 sky130_fd_sc_hd__buf_1 _10579_ (.A(_05185_),
    .X(_00041_));
 sky130_fd_sc_hd__o21a_2 _10580_ (.A1(_05085_),
    .A2(_05149_),
    .B1(net535),
    .X(_05186_));
 sky130_fd_sc_hd__a31o_2 _10581_ (.A1(_04898_),
    .A2(_05183_),
    .A3(_05146_),
    .B1(_05186_),
    .X(_00042_));
 sky130_fd_sc_hd__buf_1 _10582_ (.A(_04903_),
    .X(_05187_));
 sky130_fd_sc_hd__mux2_2 _10583_ (.A0(_05187_),
    .A1(net334),
    .S(_05151_),
    .X(_05188_));
 sky130_fd_sc_hd__buf_1 _10584_ (.A(_05188_),
    .X(_00043_));
 sky130_fd_sc_hd__inv_2 _10585_ (.A(net64),
    .Y(_05189_));
 sky130_fd_sc_hd__o21ai_2 _10586_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_05143_),
    .Y(_05190_));
 sky130_fd_sc_hd__o21ai_2 _10587_ (.A1(_05189_),
    .A2(_05143_),
    .B1(_05190_),
    .Y(_00044_));
 sky130_fd_sc_hd__and4b_2 _10588_ (.A_N(_04918_),
    .B(_04728_),
    .C(_04922_),
    .D(_04916_),
    .X(_05191_));
 sky130_fd_sc_hd__nor2_2 _10589_ (.A(net34),
    .B(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__a21oi_2 _10590_ (.A1(_04719_),
    .A2(_05191_),
    .B1(_05192_),
    .Y(_00045_));
 sky130_fd_sc_hd__nand4b_2 _10591_ (.A_N(_04917_),
    .B(_04727_),
    .C(_04922_),
    .D(_04915_),
    .Y(_05193_));
 sky130_fd_sc_hd__buf_1 _10592_ (.A(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__mux2_2 _10593_ (.A0(_04736_),
    .A1(net735),
    .S(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__buf_1 _10594_ (.A(_05195_),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_2 _10595_ (.A0(_04747_),
    .A1(\rvsingle.dp.rf.rf[22][2] ),
    .S(_05194_),
    .X(_05196_));
 sky130_fd_sc_hd__buf_1 _10596_ (.A(_05196_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_2 _10597_ (.A0(_04755_),
    .A1(net802),
    .S(_05194_),
    .X(_05197_));
 sky130_fd_sc_hd__buf_1 _10598_ (.A(_05197_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_2 _10599_ (.A0(_04760_),
    .A1(net672),
    .S(_05194_),
    .X(_05198_));
 sky130_fd_sc_hd__buf_1 _10600_ (.A(_05198_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_2 _10601_ (.A0(_04765_),
    .A1(\rvsingle.dp.rf.rf[22][5] ),
    .S(_05194_),
    .X(_05199_));
 sky130_fd_sc_hd__buf_1 _10602_ (.A(_05199_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_2 _10603_ (.A0(_04770_),
    .A1(\rvsingle.dp.rf.rf[22][6] ),
    .S(_05194_),
    .X(_05200_));
 sky130_fd_sc_hd__buf_1 _10604_ (.A(_05200_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_2 _10605_ (.A0(_04774_),
    .A1(net575),
    .S(_05194_),
    .X(_05201_));
 sky130_fd_sc_hd__buf_1 _10606_ (.A(_05201_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_2 _10607_ (.A0(_04778_),
    .A1(\rvsingle.dp.rf.rf[22][8] ),
    .S(_05194_),
    .X(_05202_));
 sky130_fd_sc_hd__buf_1 _10608_ (.A(_05202_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_2 _10609_ (.A0(_04782_),
    .A1(net479),
    .S(_05194_),
    .X(_05203_));
 sky130_fd_sc_hd__buf_1 _10610_ (.A(_05203_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_2 _10611_ (.A0(_04786_),
    .A1(net694),
    .S(_05194_),
    .X(_05204_));
 sky130_fd_sc_hd__buf_1 _10612_ (.A(_05204_),
    .X(_00055_));
 sky130_fd_sc_hd__buf_1 _10613_ (.A(_05193_),
    .X(_05205_));
 sky130_fd_sc_hd__mux2_2 _10614_ (.A0(_04790_),
    .A1(net745),
    .S(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__buf_1 _10615_ (.A(_05206_),
    .X(_00056_));
 sky130_fd_sc_hd__buf_1 _10616_ (.A(_04794_),
    .X(_05207_));
 sky130_fd_sc_hd__mux2_2 _10617_ (.A0(_05207_),
    .A1(\rvsingle.dp.rf.rf[22][12] ),
    .S(_05205_),
    .X(_05208_));
 sky130_fd_sc_hd__buf_1 _10618_ (.A(_05208_),
    .X(_00057_));
 sky130_fd_sc_hd__buf_1 _10619_ (.A(_04800_),
    .X(_05209_));
 sky130_fd_sc_hd__mux2_2 _10620_ (.A0(_05209_),
    .A1(\rvsingle.dp.rf.rf[22][13] ),
    .S(_05205_),
    .X(_05210_));
 sky130_fd_sc_hd__buf_1 _10621_ (.A(_05210_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_2 _10622_ (.A0(_04808_),
    .A1(\rvsingle.dp.rf.rf[22][14] ),
    .S(_05205_),
    .X(_05211_));
 sky130_fd_sc_hd__buf_1 _10623_ (.A(_05211_),
    .X(_00059_));
 sky130_fd_sc_hd__buf_1 _10624_ (.A(_04813_),
    .X(_05212_));
 sky130_fd_sc_hd__mux2_2 _10625_ (.A0(_05212_),
    .A1(\rvsingle.dp.rf.rf[22][15] ),
    .S(_05205_),
    .X(_05213_));
 sky130_fd_sc_hd__buf_1 _10626_ (.A(_05213_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_2 _10627_ (.A0(_04818_),
    .A1(net711),
    .S(_05205_),
    .X(_05214_));
 sky130_fd_sc_hd__buf_1 _10628_ (.A(_05214_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_2 _10629_ (.A0(_04824_),
    .A1(net369),
    .S(_05205_),
    .X(_05215_));
 sky130_fd_sc_hd__buf_1 _10630_ (.A(_05215_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_2 _10631_ (.A0(_04828_),
    .A1(net558),
    .S(_05205_),
    .X(_05216_));
 sky130_fd_sc_hd__buf_1 _10632_ (.A(_05216_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_2 _10633_ (.A0(_04834_),
    .A1(net507),
    .S(_05205_),
    .X(_05217_));
 sky130_fd_sc_hd__buf_1 _10634_ (.A(_05217_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_2 _10635_ (.A0(_04840_),
    .A1(net609),
    .S(_05205_),
    .X(_05218_));
 sky130_fd_sc_hd__buf_1 _10636_ (.A(_05218_),
    .X(_00065_));
 sky130_fd_sc_hd__buf_1 _10637_ (.A(_05193_),
    .X(_05219_));
 sky130_fd_sc_hd__mux2_2 _10638_ (.A0(_04846_),
    .A1(net347),
    .S(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__buf_1 _10639_ (.A(_05220_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_2 _10640_ (.A0(_04853_),
    .A1(net754),
    .S(_05219_),
    .X(_05221_));
 sky130_fd_sc_hd__buf_1 _10641_ (.A(_05221_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_2 _10642_ (.A0(_04859_),
    .A1(net567),
    .S(_05219_),
    .X(_05222_));
 sky130_fd_sc_hd__buf_1 _10643_ (.A(_05222_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_2 _10644_ (.A0(_04863_),
    .A1(net514),
    .S(_05219_),
    .X(_05223_));
 sky130_fd_sc_hd__buf_1 _10645_ (.A(_05223_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_2 _10646_ (.A0(_04870_),
    .A1(net747),
    .S(_05219_),
    .X(_05224_));
 sky130_fd_sc_hd__buf_1 _10647_ (.A(_05224_),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_2 _10648_ (.A0(_04877_),
    .A1(net546),
    .S(_05219_),
    .X(_05225_));
 sky130_fd_sc_hd__buf_1 _10649_ (.A(_05225_),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_2 _10650_ (.A0(_04886_),
    .A1(net662),
    .S(_05219_),
    .X(_05226_));
 sky130_fd_sc_hd__buf_1 _10651_ (.A(_05226_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_2 _10652_ (.A0(_04892_),
    .A1(net330),
    .S(_05219_),
    .X(_05227_));
 sky130_fd_sc_hd__buf_1 _10653_ (.A(_05227_),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_2 _10654_ (.A0(_04898_),
    .A1(net624),
    .S(_05219_),
    .X(_05228_));
 sky130_fd_sc_hd__buf_1 _10655_ (.A(_05228_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_2 _10656_ (.A0(_05187_),
    .A1(net402),
    .S(_05219_),
    .X(_05229_));
 sky130_fd_sc_hd__buf_1 _10657_ (.A(_05229_),
    .X(_00075_));
 sky130_fd_sc_hd__inv_2 _10658_ (.A(net40),
    .Y(_05230_));
 sky130_fd_sc_hd__o21ai_2 _10659_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_05191_),
    .Y(_05231_));
 sky130_fd_sc_hd__o21ai_2 _10660_ (.A1(_05230_),
    .A2(_05191_),
    .B1(_05231_),
    .Y(_00076_));
 sky130_fd_sc_hd__and4b_2 _10661_ (.A_N(_04918_),
    .B(_04922_),
    .C(_05057_),
    .D(_04916_),
    .X(_05232_));
 sky130_fd_sc_hd__nor2_2 _10662_ (.A(net127),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__a21oi_2 _10663_ (.A1(_04719_),
    .A2(_05232_),
    .B1(_05233_),
    .Y(_00077_));
 sky130_fd_sc_hd__or4bb_2 _10664_ (.A(_04917_),
    .B(_04928_),
    .C_N(_05057_),
    .D_N(_04915_),
    .X(_05234_));
 sky130_fd_sc_hd__buf_1 _10665_ (.A(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__mux2_2 _10666_ (.A0(_04736_),
    .A1(net499),
    .S(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__buf_1 _10667_ (.A(_05236_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_2 _10668_ (.A0(_04747_),
    .A1(net783),
    .S(_05235_),
    .X(_05237_));
 sky130_fd_sc_hd__buf_1 _10669_ (.A(_05237_),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_2 _10670_ (.A0(_04755_),
    .A1(net454),
    .S(_05235_),
    .X(_05238_));
 sky130_fd_sc_hd__buf_1 _10671_ (.A(_05238_),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_2 _10672_ (.A0(_04760_),
    .A1(\rvsingle.dp.rf.rf[21][4] ),
    .S(_05235_),
    .X(_05239_));
 sky130_fd_sc_hd__buf_1 _10673_ (.A(_05239_),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_2 _10674_ (.A0(_04765_),
    .A1(net650),
    .S(_05235_),
    .X(_05240_));
 sky130_fd_sc_hd__buf_1 _10675_ (.A(_05240_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_2 _10676_ (.A0(_04770_),
    .A1(\rvsingle.dp.rf.rf[21][6] ),
    .S(_05235_),
    .X(_05241_));
 sky130_fd_sc_hd__buf_1 _10677_ (.A(_05241_),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_2 _10678_ (.A0(_04774_),
    .A1(net318),
    .S(_05235_),
    .X(_05242_));
 sky130_fd_sc_hd__buf_1 _10679_ (.A(_05242_),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_2 _10680_ (.A0(_04778_),
    .A1(net683),
    .S(_05235_),
    .X(_05243_));
 sky130_fd_sc_hd__buf_1 _10681_ (.A(_05243_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_2 _10682_ (.A0(_04782_),
    .A1(net325),
    .S(_05235_),
    .X(_05244_));
 sky130_fd_sc_hd__buf_1 _10683_ (.A(_05244_),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_2 _10684_ (.A0(_04786_),
    .A1(\rvsingle.dp.rf.rf[21][10] ),
    .S(_05235_),
    .X(_05245_));
 sky130_fd_sc_hd__buf_1 _10685_ (.A(_05245_),
    .X(_00087_));
 sky130_fd_sc_hd__buf_1 _10686_ (.A(_05234_),
    .X(_05246_));
 sky130_fd_sc_hd__mux2_2 _10687_ (.A0(_04790_),
    .A1(\rvsingle.dp.rf.rf[21][11] ),
    .S(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__buf_1 _10688_ (.A(_05247_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_2 _10689_ (.A0(_05207_),
    .A1(net423),
    .S(_05246_),
    .X(_05248_));
 sky130_fd_sc_hd__buf_1 _10690_ (.A(_05248_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_2 _10691_ (.A0(_05209_),
    .A1(\rvsingle.dp.rf.rf[21][13] ),
    .S(_05246_),
    .X(_05249_));
 sky130_fd_sc_hd__buf_1 _10692_ (.A(_05249_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_2 _10693_ (.A0(_04808_),
    .A1(\rvsingle.dp.rf.rf[21][14] ),
    .S(_05246_),
    .X(_05250_));
 sky130_fd_sc_hd__buf_1 _10694_ (.A(_05250_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_2 _10695_ (.A0(_05212_),
    .A1(net500),
    .S(_05246_),
    .X(_05251_));
 sky130_fd_sc_hd__buf_1 _10696_ (.A(_05251_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_2 _10697_ (.A0(_04818_),
    .A1(net345),
    .S(_05246_),
    .X(_05252_));
 sky130_fd_sc_hd__buf_1 _10698_ (.A(_05252_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_2 _10699_ (.A0(_04824_),
    .A1(net630),
    .S(_05246_),
    .X(_05253_));
 sky130_fd_sc_hd__buf_1 _10700_ (.A(_05253_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_2 _10701_ (.A0(_04828_),
    .A1(net521),
    .S(_05246_),
    .X(_05254_));
 sky130_fd_sc_hd__buf_1 _10702_ (.A(_05254_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_2 _10703_ (.A0(_04834_),
    .A1(\rvsingle.dp.rf.rf[21][19] ),
    .S(_05246_),
    .X(_05255_));
 sky130_fd_sc_hd__buf_1 _10704_ (.A(_05255_),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_2 _10705_ (.A0(_04840_),
    .A1(net548),
    .S(_05246_),
    .X(_05256_));
 sky130_fd_sc_hd__buf_1 _10706_ (.A(_05256_),
    .X(_00097_));
 sky130_fd_sc_hd__buf_1 _10707_ (.A(_05234_),
    .X(_05257_));
 sky130_fd_sc_hd__mux2_2 _10708_ (.A0(_04846_),
    .A1(\rvsingle.dp.rf.rf[21][21] ),
    .S(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__buf_1 _10709_ (.A(_05258_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_2 _10710_ (.A0(_04853_),
    .A1(net670),
    .S(_05257_),
    .X(_05259_));
 sky130_fd_sc_hd__buf_1 _10711_ (.A(_05259_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_2 _10712_ (.A0(_04859_),
    .A1(net619),
    .S(_05257_),
    .X(_05260_));
 sky130_fd_sc_hd__buf_1 _10713_ (.A(_05260_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_2 _10714_ (.A0(_04863_),
    .A1(net411),
    .S(_05257_),
    .X(_05261_));
 sky130_fd_sc_hd__buf_1 _10715_ (.A(_05261_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_2 _10716_ (.A0(_04870_),
    .A1(net365),
    .S(_05257_),
    .X(_05262_));
 sky130_fd_sc_hd__buf_1 _10717_ (.A(_05262_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_2 _10718_ (.A0(_04877_),
    .A1(net756),
    .S(_05257_),
    .X(_05263_));
 sky130_fd_sc_hd__buf_1 _10719_ (.A(_05263_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_2 _10720_ (.A0(_04886_),
    .A1(net750),
    .S(_05257_),
    .X(_05264_));
 sky130_fd_sc_hd__buf_1 _10721_ (.A(_05264_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_2 _10722_ (.A0(_04892_),
    .A1(net430),
    .S(_05257_),
    .X(_05265_));
 sky130_fd_sc_hd__buf_1 _10723_ (.A(_05265_),
    .X(_00105_));
 sky130_fd_sc_hd__buf_1 _10724_ (.A(_04897_),
    .X(_05266_));
 sky130_fd_sc_hd__mux2_2 _10725_ (.A0(_05266_),
    .A1(net773),
    .S(_05257_),
    .X(_05267_));
 sky130_fd_sc_hd__buf_1 _10726_ (.A(_05267_),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_2 _10727_ (.A0(_05187_),
    .A1(net326),
    .S(_05257_),
    .X(_05268_));
 sky130_fd_sc_hd__buf_1 _10728_ (.A(_05268_),
    .X(_00107_));
 sky130_fd_sc_hd__inv_2 _10729_ (.A(net58),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_2 _10730_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_05232_),
    .Y(_05270_));
 sky130_fd_sc_hd__o21ai_2 _10731_ (.A1(_05269_),
    .A2(_05232_),
    .B1(_05270_),
    .Y(_00108_));
 sky130_fd_sc_hd__and4b_2 _10732_ (.A_N(_04917_),
    .B(_04920_),
    .C(_04922_),
    .D(_04916_),
    .X(_05271_));
 sky130_fd_sc_hd__nor2_2 _10733_ (.A(net9),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__a21oi_2 _10734_ (.A1(_04719_),
    .A2(_05271_),
    .B1(_05272_),
    .Y(_00109_));
 sky130_fd_sc_hd__nand4b_2 _10735_ (.A_N(_04917_),
    .B(_04920_),
    .C(_04921_),
    .D(_04915_),
    .Y(_05273_));
 sky130_fd_sc_hd__buf_1 _10736_ (.A(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__mux2_2 _10737_ (.A0(_04736_),
    .A1(\rvsingle.dp.rf.rf[20][1] ),
    .S(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__buf_1 _10738_ (.A(_05275_),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_2 _10739_ (.A0(_04747_),
    .A1(net790),
    .S(_05274_),
    .X(_05276_));
 sky130_fd_sc_hd__buf_1 _10740_ (.A(_05276_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_2 _10741_ (.A0(_04755_),
    .A1(\rvsingle.dp.rf.rf[20][3] ),
    .S(_05274_),
    .X(_05277_));
 sky130_fd_sc_hd__buf_1 _10742_ (.A(_05277_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_2 _10743_ (.A0(_04760_),
    .A1(net807),
    .S(_05274_),
    .X(_05278_));
 sky130_fd_sc_hd__buf_1 _10744_ (.A(_05278_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_2 _10745_ (.A0(_04765_),
    .A1(\rvsingle.dp.rf.rf[20][5] ),
    .S(_05274_),
    .X(_05279_));
 sky130_fd_sc_hd__buf_1 _10746_ (.A(_05279_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_2 _10747_ (.A0(_04770_),
    .A1(\rvsingle.dp.rf.rf[20][6] ),
    .S(_05274_),
    .X(_05280_));
 sky130_fd_sc_hd__buf_1 _10748_ (.A(_05280_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_2 _10749_ (.A0(_04774_),
    .A1(\rvsingle.dp.rf.rf[20][7] ),
    .S(_05274_),
    .X(_05281_));
 sky130_fd_sc_hd__buf_1 _10750_ (.A(_05281_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_2 _10751_ (.A0(_04778_),
    .A1(\rvsingle.dp.rf.rf[20][8] ),
    .S(_05274_),
    .X(_05282_));
 sky130_fd_sc_hd__buf_1 _10752_ (.A(_05282_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_2 _10753_ (.A0(_04782_),
    .A1(net583),
    .S(_05274_),
    .X(_05283_));
 sky130_fd_sc_hd__buf_1 _10754_ (.A(_05283_),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_2 _10755_ (.A0(_04786_),
    .A1(net782),
    .S(_05274_),
    .X(_05284_));
 sky130_fd_sc_hd__buf_1 _10756_ (.A(_05284_),
    .X(_00119_));
 sky130_fd_sc_hd__buf_1 _10757_ (.A(_05273_),
    .X(_05285_));
 sky130_fd_sc_hd__mux2_2 _10758_ (.A0(_04790_),
    .A1(\rvsingle.dp.rf.rf[20][11] ),
    .S(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__buf_1 _10759_ (.A(_05286_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_2 _10760_ (.A0(_05207_),
    .A1(\rvsingle.dp.rf.rf[20][12] ),
    .S(_05285_),
    .X(_05287_));
 sky130_fd_sc_hd__buf_1 _10761_ (.A(_05287_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_2 _10762_ (.A0(_05209_),
    .A1(\rvsingle.dp.rf.rf[20][13] ),
    .S(_05285_),
    .X(_05288_));
 sky130_fd_sc_hd__buf_1 _10763_ (.A(_05288_),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_2 _10764_ (.A0(_04808_),
    .A1(net647),
    .S(_05285_),
    .X(_05289_));
 sky130_fd_sc_hd__buf_1 _10765_ (.A(_05289_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_2 _10766_ (.A0(_05212_),
    .A1(\rvsingle.dp.rf.rf[20][15] ),
    .S(_05285_),
    .X(_05290_));
 sky130_fd_sc_hd__buf_1 _10767_ (.A(_05290_),
    .X(_00124_));
 sky130_fd_sc_hd__buf_1 _10768_ (.A(_04817_),
    .X(_05291_));
 sky130_fd_sc_hd__mux2_2 _10769_ (.A0(_05291_),
    .A1(net739),
    .S(_05285_),
    .X(_05292_));
 sky130_fd_sc_hd__buf_1 _10770_ (.A(_05292_),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_2 _10771_ (.A0(_04824_),
    .A1(net485),
    .S(_05285_),
    .X(_05293_));
 sky130_fd_sc_hd__buf_1 _10772_ (.A(_05293_),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_2 _10773_ (.A0(_04828_),
    .A1(\rvsingle.dp.rf.rf[20][18] ),
    .S(_05285_),
    .X(_05294_));
 sky130_fd_sc_hd__buf_1 _10774_ (.A(_05294_),
    .X(_00127_));
 sky130_fd_sc_hd__buf_1 _10775_ (.A(_04833_),
    .X(_05295_));
 sky130_fd_sc_hd__mux2_2 _10776_ (.A0(_05295_),
    .A1(net685),
    .S(_05285_),
    .X(_05296_));
 sky130_fd_sc_hd__buf_1 _10777_ (.A(_05296_),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_2 _10778_ (.A0(_04840_),
    .A1(net794),
    .S(_05285_),
    .X(_05297_));
 sky130_fd_sc_hd__buf_1 _10779_ (.A(_05297_),
    .X(_00129_));
 sky130_fd_sc_hd__buf_1 _10780_ (.A(_05273_),
    .X(_05298_));
 sky130_fd_sc_hd__mux2_2 _10781_ (.A0(_04846_),
    .A1(net571),
    .S(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__buf_1 _10782_ (.A(_05299_),
    .X(_00130_));
 sky130_fd_sc_hd__buf_1 _10783_ (.A(_04852_),
    .X(_05300_));
 sky130_fd_sc_hd__mux2_2 _10784_ (.A0(_05300_),
    .A1(net463),
    .S(_05298_),
    .X(_05301_));
 sky130_fd_sc_hd__buf_1 _10785_ (.A(_05301_),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_2 _10786_ (.A0(_04859_),
    .A1(net424),
    .S(_05298_),
    .X(_05302_));
 sky130_fd_sc_hd__buf_1 _10787_ (.A(_05302_),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_2 _10788_ (.A0(_04863_),
    .A1(net413),
    .S(_05298_),
    .X(_05303_));
 sky130_fd_sc_hd__buf_1 _10789_ (.A(_05303_),
    .X(_00133_));
 sky130_fd_sc_hd__buf_1 _10790_ (.A(_04868_),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_2 _10791_ (.A0(_05304_),
    .A1(net589),
    .S(_05298_),
    .X(_05305_));
 sky130_fd_sc_hd__buf_1 _10792_ (.A(_05305_),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_2 _10793_ (.A0(_04877_),
    .A1(net591),
    .S(_05298_),
    .X(_05306_));
 sky130_fd_sc_hd__buf_1 _10794_ (.A(_05306_),
    .X(_00135_));
 sky130_fd_sc_hd__buf_1 _10795_ (.A(_04885_),
    .X(_05307_));
 sky130_fd_sc_hd__mux2_2 _10796_ (.A0(_05307_),
    .A1(net517),
    .S(_05298_),
    .X(_05308_));
 sky130_fd_sc_hd__buf_1 _10797_ (.A(_05308_),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_2 _10798_ (.A0(_04892_),
    .A1(net344),
    .S(_05298_),
    .X(_05309_));
 sky130_fd_sc_hd__buf_1 _10799_ (.A(_05309_),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_2 _10800_ (.A0(_05266_),
    .A1(net461),
    .S(_05298_),
    .X(_05310_));
 sky130_fd_sc_hd__buf_1 _10801_ (.A(_05310_),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_2 _10802_ (.A0(_05187_),
    .A1(net447),
    .S(_05298_),
    .X(_05311_));
 sky130_fd_sc_hd__buf_1 _10803_ (.A(_05311_),
    .X(_00139_));
 sky130_fd_sc_hd__inv_2 _10804_ (.A(net47),
    .Y(_05312_));
 sky130_fd_sc_hd__o21ai_2 _10805_ (.A1(_04909_),
    .A2(_04913_),
    .B1(_05271_),
    .Y(_05313_));
 sky130_fd_sc_hd__o21ai_2 _10806_ (.A1(_05312_),
    .A2(_05271_),
    .B1(_05313_),
    .Y(_00140_));
 sky130_fd_sc_hd__buf_1 _10807_ (.A(_04718_),
    .X(_05314_));
 sky130_fd_sc_hd__and3_2 _10808_ (.A(_05097_),
    .B(_04726_),
    .C(_05058_),
    .X(_05315_));
 sky130_fd_sc_hd__buf_1 _10809_ (.A(_04725_),
    .X(_05316_));
 sky130_fd_sc_hd__a21oi_2 _10810_ (.A1(_05316_),
    .A2(_05145_),
    .B1(net4),
    .Y(_05317_));
 sky130_fd_sc_hd__a21oi_2 _10811_ (.A1(_05314_),
    .A2(_05315_),
    .B1(_05317_),
    .Y(_00141_));
 sky130_fd_sc_hd__buf_1 _10812_ (.A(_04735_),
    .X(_05318_));
 sky130_fd_sc_hd__or4_2 _10813_ (.A(_04722_),
    .B(_04723_),
    .C(_04965_),
    .D(_05063_),
    .X(_05319_));
 sky130_fd_sc_hd__buf_1 _10814_ (.A(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_2 _10815_ (.A0(_05318_),
    .A1(net280),
    .S(_05320_),
    .X(_05321_));
 sky130_fd_sc_hd__buf_1 _10816_ (.A(_05321_),
    .X(_00142_));
 sky130_fd_sc_hd__buf_1 _10817_ (.A(_04746_),
    .X(_05322_));
 sky130_fd_sc_hd__mux2_2 _10818_ (.A0(_05322_),
    .A1(net638),
    .S(_05320_),
    .X(_05323_));
 sky130_fd_sc_hd__buf_1 _10819_ (.A(_05323_),
    .X(_00143_));
 sky130_fd_sc_hd__or4b_2 _10820_ (.A(_04982_),
    .B(_04983_),
    .C(_04981_),
    .D_N(_04754_),
    .X(_05324_));
 sky130_fd_sc_hd__buf_1 _10821_ (.A(_05320_),
    .X(_05325_));
 sky130_fd_sc_hd__a2bb2o_2 _10822_ (.A1_N(_05085_),
    .A2_N(_05324_),
    .B1(_05325_),
    .B2(net118),
    .X(_00144_));
 sky130_fd_sc_hd__or4b_2 _10823_ (.A(_04982_),
    .B(_04983_),
    .C(_04981_),
    .D_N(_04759_),
    .X(_05326_));
 sky130_fd_sc_hd__a2bb2o_2 _10824_ (.A1_N(_05085_),
    .A2_N(_05326_),
    .B1(_05325_),
    .B2(net193),
    .X(_00145_));
 sky130_fd_sc_hd__and2_2 _10825_ (.A(_04764_),
    .B(_05316_),
    .X(_05327_));
 sky130_fd_sc_hd__a32o_2 _10826_ (.A1(_05327_),
    .A2(_05069_),
    .A3(_05068_),
    .B1(_05325_),
    .B2(net13),
    .X(_00146_));
 sky130_fd_sc_hd__or4b_2 _10827_ (.A(_04982_),
    .B(_04983_),
    .C(_04981_),
    .D_N(_04769_),
    .X(_05328_));
 sky130_fd_sc_hd__a2bb2o_2 _10828_ (.A1_N(_05085_),
    .A2_N(_05328_),
    .B1(_05325_),
    .B2(net210),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_2 _10829_ (.A0(_04774_),
    .A1(net383),
    .S(_05320_),
    .X(_05329_));
 sky130_fd_sc_hd__buf_1 _10830_ (.A(_05329_),
    .X(_00148_));
 sky130_fd_sc_hd__buf_1 _10831_ (.A(_04777_),
    .X(_05330_));
 sky130_fd_sc_hd__mux2_2 _10832_ (.A0(_05330_),
    .A1(net704),
    .S(_05320_),
    .X(_05331_));
 sky130_fd_sc_hd__buf_1 _10833_ (.A(_05331_),
    .X(_00149_));
 sky130_fd_sc_hd__and2_2 _10834_ (.A(_04781_),
    .B(_04726_),
    .X(_05332_));
 sky130_fd_sc_hd__a32o_2 _10835_ (.A1(_05332_),
    .A2(_05069_),
    .A3(_05068_),
    .B1(_05325_),
    .B2(net3),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_2 _10836_ (.A0(_04786_),
    .A1(net489),
    .S(_05320_),
    .X(_05333_));
 sky130_fd_sc_hd__buf_1 _10837_ (.A(_05333_),
    .X(_00151_));
 sky130_fd_sc_hd__buf_1 _10838_ (.A(_04789_),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_2 _10839_ (.A0(_05334_),
    .A1(net342),
    .S(_05320_),
    .X(_05335_));
 sky130_fd_sc_hd__buf_1 _10840_ (.A(_05335_),
    .X(_00152_));
 sky130_fd_sc_hd__buf_1 _10841_ (.A(_05316_),
    .X(_05336_));
 sky130_fd_sc_hd__buf_1 _10842_ (.A(_04915_),
    .X(_05337_));
 sky130_fd_sc_hd__buf_1 _10843_ (.A(_04917_),
    .X(_05338_));
 sky130_fd_sc_hd__buf_1 _10844_ (.A(_04965_),
    .X(_05339_));
 sky130_fd_sc_hd__o41a_2 _10845_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05084_),
    .B1(net184),
    .X(_05340_));
 sky130_fd_sc_hd__a31o_2 _10846_ (.A1(_04796_),
    .A2(_05183_),
    .A3(_05336_),
    .B1(_05340_),
    .X(_00153_));
 sky130_fd_sc_hd__o41a_2 _10847_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05084_),
    .B1(net195),
    .X(_05341_));
 sky130_fd_sc_hd__a31o_2 _10848_ (.A1(_04802_),
    .A2(_05183_),
    .A3(_05336_),
    .B1(_05341_),
    .X(_00154_));
 sky130_fd_sc_hd__or4b_2 _10849_ (.A(_04916_),
    .B(_04918_),
    .C(_04965_),
    .D_N(_04807_),
    .X(_05342_));
 sky130_fd_sc_hd__a2bb2o_2 _10850_ (.A1_N(_05085_),
    .A2_N(_05342_),
    .B1(_05325_),
    .B2(net98),
    .X(_00155_));
 sky130_fd_sc_hd__nand2_2 _10851_ (.A(_04814_),
    .B(_05316_),
    .Y(_05343_));
 sky130_fd_sc_hd__a2bb2o_2 _10852_ (.A1_N(_05085_),
    .A2_N(_05343_),
    .B1(_05325_),
    .B2(net132),
    .X(_00156_));
 sky130_fd_sc_hd__buf_1 _10853_ (.A(_04817_),
    .X(_05344_));
 sky130_fd_sc_hd__and2_2 _10854_ (.A(_05344_),
    .B(_04726_),
    .X(_05345_));
 sky130_fd_sc_hd__a32o_2 _10855_ (.A1(_05345_),
    .A2(_05069_),
    .A3(_05068_),
    .B1(_05325_),
    .B2(net22),
    .X(_00157_));
 sky130_fd_sc_hd__and2_2 _10856_ (.A(_04823_),
    .B(_04726_),
    .X(_05346_));
 sky130_fd_sc_hd__a32o_2 _10857_ (.A1(_05346_),
    .A2(_05069_),
    .A3(_05068_),
    .B1(_05320_),
    .B2(net39),
    .X(_00158_));
 sky130_fd_sc_hd__and2_2 _10858_ (.A(_05173_),
    .B(_04726_),
    .X(_05347_));
 sky130_fd_sc_hd__a32o_2 _10859_ (.A1(_05347_),
    .A2(_05069_),
    .A3(_05068_),
    .B1(_05320_),
    .B2(net12),
    .X(_00159_));
 sky130_fd_sc_hd__nand2_2 _10860_ (.A(_04834_),
    .B(_05316_),
    .Y(_05348_));
 sky130_fd_sc_hd__a2bb2o_2 _10861_ (.A1_N(_05085_),
    .A2_N(_05348_),
    .B1(_05325_),
    .B2(net169),
    .X(_00160_));
 sky130_fd_sc_hd__o41a_2 _10862_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05084_),
    .B1(net205),
    .X(_05349_));
 sky130_fd_sc_hd__a31o_2 _10863_ (.A1(_04840_),
    .A2(_05183_),
    .A3(_05336_),
    .B1(_05349_),
    .X(_00161_));
 sky130_fd_sc_hd__nand2_2 _10864_ (.A(_04846_),
    .B(_05316_),
    .Y(_05350_));
 sky130_fd_sc_hd__a2bb2o_2 _10865_ (.A1_N(_05085_),
    .A2_N(_05350_),
    .B1(_05325_),
    .B2(net145),
    .X(_00162_));
 sky130_fd_sc_hd__o41a_2 _10866_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05084_),
    .B1(net206),
    .X(_05351_));
 sky130_fd_sc_hd__a31o_2 _10867_ (.A1(_04853_),
    .A2(_05183_),
    .A3(_05336_),
    .B1(_05351_),
    .X(_00163_));
 sky130_fd_sc_hd__buf_1 _10868_ (.A(_04858_),
    .X(_05352_));
 sky130_fd_sc_hd__mux2_2 _10869_ (.A0(_05352_),
    .A1(net238),
    .S(_05320_),
    .X(_05353_));
 sky130_fd_sc_hd__buf_1 _10870_ (.A(_05353_),
    .X(_00164_));
 sky130_fd_sc_hd__buf_1 _10871_ (.A(_04862_),
    .X(_05354_));
 sky130_fd_sc_hd__mux2_2 _10872_ (.A0(_05354_),
    .A1(net244),
    .S(_05319_),
    .X(_05355_));
 sky130_fd_sc_hd__buf_1 _10873_ (.A(_05355_),
    .X(_00165_));
 sky130_fd_sc_hd__o41a_2 _10874_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05084_),
    .B1(net319),
    .X(_05356_));
 sky130_fd_sc_hd__a31o_2 _10875_ (.A1(_04870_),
    .A2(_05183_),
    .A3(_05336_),
    .B1(_05356_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_2 _10876_ (.A0(_04877_),
    .A1(net296),
    .S(_05319_),
    .X(_05357_));
 sky130_fd_sc_hd__buf_1 _10877_ (.A(_05357_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_2 _10878_ (.A0(_05307_),
    .A1(\rvsingle.dp.rf.rf[1][27] ),
    .S(_05319_),
    .X(_05358_));
 sky130_fd_sc_hd__buf_1 _10879_ (.A(_05358_),
    .X(_00168_));
 sky130_fd_sc_hd__buf_1 _10880_ (.A(_04891_),
    .X(_05359_));
 sky130_fd_sc_hd__mux2_2 _10881_ (.A0(_05359_),
    .A1(net641),
    .S(_05319_),
    .X(_05360_));
 sky130_fd_sc_hd__buf_1 _10882_ (.A(_05360_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_2 _10883_ (.A0(_05266_),
    .A1(\rvsingle.dp.rf.rf[1][29] ),
    .S(_05319_),
    .X(_05361_));
 sky130_fd_sc_hd__buf_1 _10884_ (.A(_05361_),
    .X(_00170_));
 sky130_fd_sc_hd__o41a_2 _10885_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05084_),
    .B1(net300),
    .X(_05362_));
 sky130_fd_sc_hd__a31o_2 _10886_ (.A1(_04904_),
    .A2(_05183_),
    .A3(_05336_),
    .B1(_05362_),
    .X(_00171_));
 sky130_fd_sc_hd__inv_2 _10887_ (.A(net73),
    .Y(_05363_));
 sky130_fd_sc_hd__buf_1 _10888_ (.A(_04908_),
    .X(_05364_));
 sky130_fd_sc_hd__buf_1 _10889_ (.A(_04912_),
    .X(_05365_));
 sky130_fd_sc_hd__o21ai_2 _10890_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05315_),
    .Y(_05366_));
 sky130_fd_sc_hd__o21ai_2 _10891_ (.A1(_05363_),
    .A2(_05315_),
    .B1(_05366_),
    .Y(_00172_));
 sky130_fd_sc_hd__nor3b_2 _10892_ (.A(_04917_),
    .B(_04965_),
    .C_N(_04915_),
    .Y(_05367_));
 sky130_fd_sc_hd__and3_2 _10893_ (.A(_04721_),
    .B(_04728_),
    .C(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__nor2_2 _10894_ (.A(net115),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__a21oi_2 _10895_ (.A1(_05314_),
    .A2(_05368_),
    .B1(_05369_),
    .Y(_00173_));
 sky130_fd_sc_hd__or3b_2 _10896_ (.A(_04723_),
    .B(_04724_),
    .C_N(_04722_),
    .X(_05370_));
 sky130_fd_sc_hd__buf_1 _10897_ (.A(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__or4b_2 _10898_ (.A(_04738_),
    .B(_04733_),
    .C(_05371_),
    .D_N(_04739_),
    .X(_05372_));
 sky130_fd_sc_hd__buf_1 _10899_ (.A(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__mux2_2 _10900_ (.A0(_05318_),
    .A1(\rvsingle.dp.rf.rf[18][1] ),
    .S(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__buf_1 _10901_ (.A(_05374_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_2 _10902_ (.A0(_05322_),
    .A1(\rvsingle.dp.rf.rf[18][2] ),
    .S(_05373_),
    .X(_05375_));
 sky130_fd_sc_hd__buf_1 _10903_ (.A(_05375_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_2 _10904_ (.A0(_04755_),
    .A1(\rvsingle.dp.rf.rf[18][3] ),
    .S(_05373_),
    .X(_05376_));
 sky130_fd_sc_hd__buf_1 _10905_ (.A(_05376_),
    .X(_00176_));
 sky130_fd_sc_hd__buf_1 _10906_ (.A(_04759_),
    .X(_05377_));
 sky130_fd_sc_hd__mux2_2 _10907_ (.A0(_05377_),
    .A1(net529),
    .S(_05373_),
    .X(_05378_));
 sky130_fd_sc_hd__buf_1 _10908_ (.A(_05378_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_2 _10909_ (.A0(_04765_),
    .A1(\rvsingle.dp.rf.rf[18][5] ),
    .S(_05373_),
    .X(_05379_));
 sky130_fd_sc_hd__buf_1 _10910_ (.A(_05379_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_2 _10911_ (.A0(_04770_),
    .A1(\rvsingle.dp.rf.rf[18][6] ),
    .S(_05373_),
    .X(_05380_));
 sky130_fd_sc_hd__buf_1 _10912_ (.A(_05380_),
    .X(_00179_));
 sky130_fd_sc_hd__buf_1 _10913_ (.A(_04773_),
    .X(_05381_));
 sky130_fd_sc_hd__mux2_2 _10914_ (.A0(_05381_),
    .A1(net491),
    .S(_05373_),
    .X(_05382_));
 sky130_fd_sc_hd__buf_1 _10915_ (.A(_05382_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_2 _10916_ (.A0(_05330_),
    .A1(net555),
    .S(_05373_),
    .X(_05383_));
 sky130_fd_sc_hd__buf_1 _10917_ (.A(_05383_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_2 _10918_ (.A0(_04782_),
    .A1(net577),
    .S(_05373_),
    .X(_05384_));
 sky130_fd_sc_hd__buf_1 _10919_ (.A(_05384_),
    .X(_00182_));
 sky130_fd_sc_hd__buf_1 _10920_ (.A(_04785_),
    .X(_05385_));
 sky130_fd_sc_hd__mux2_2 _10921_ (.A0(_05385_),
    .A1(net557),
    .S(_05373_),
    .X(_05386_));
 sky130_fd_sc_hd__buf_1 _10922_ (.A(_05386_),
    .X(_00183_));
 sky130_fd_sc_hd__buf_1 _10923_ (.A(_05372_),
    .X(_05387_));
 sky130_fd_sc_hd__mux2_2 _10924_ (.A0(_05334_),
    .A1(net712),
    .S(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__buf_1 _10925_ (.A(_05388_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_2 _10926_ (.A0(_05207_),
    .A1(\rvsingle.dp.rf.rf[18][12] ),
    .S(_05387_),
    .X(_05389_));
 sky130_fd_sc_hd__buf_1 _10927_ (.A(_05389_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_2 _10928_ (.A0(_05209_),
    .A1(net817),
    .S(_05387_),
    .X(_05390_));
 sky130_fd_sc_hd__buf_1 _10929_ (.A(_05390_),
    .X(_00186_));
 sky130_fd_sc_hd__buf_1 _10930_ (.A(_04807_),
    .X(_05391_));
 sky130_fd_sc_hd__mux2_2 _10931_ (.A0(_05391_),
    .A1(\rvsingle.dp.rf.rf[18][14] ),
    .S(_05387_),
    .X(_05392_));
 sky130_fd_sc_hd__buf_1 _10932_ (.A(_05392_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_2 _10933_ (.A0(_05212_),
    .A1(\rvsingle.dp.rf.rf[18][15] ),
    .S(_05387_),
    .X(_05393_));
 sky130_fd_sc_hd__buf_1 _10934_ (.A(_05393_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_2 _10935_ (.A0(_05291_),
    .A1(\rvsingle.dp.rf.rf[18][16] ),
    .S(_05387_),
    .X(_05394_));
 sky130_fd_sc_hd__buf_1 _10936_ (.A(_05394_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_2 _10937_ (.A0(_04824_),
    .A1(net349),
    .S(_05387_),
    .X(_05395_));
 sky130_fd_sc_hd__buf_1 _10938_ (.A(_05395_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_2 _10939_ (.A0(_04828_),
    .A1(net614),
    .S(_05387_),
    .X(_05396_));
 sky130_fd_sc_hd__buf_1 _10940_ (.A(_05396_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_2 _10941_ (.A0(_05295_),
    .A1(\rvsingle.dp.rf.rf[18][19] ),
    .S(_05387_),
    .X(_05397_));
 sky130_fd_sc_hd__buf_1 _10942_ (.A(_05397_),
    .X(_00192_));
 sky130_fd_sc_hd__buf_1 _10943_ (.A(_04839_),
    .X(_05398_));
 sky130_fd_sc_hd__mux2_2 _10944_ (.A0(_05398_),
    .A1(\rvsingle.dp.rf.rf[18][20] ),
    .S(_05387_),
    .X(_05399_));
 sky130_fd_sc_hd__buf_1 _10945_ (.A(_05399_),
    .X(_00193_));
 sky130_fd_sc_hd__buf_1 _10946_ (.A(_04845_),
    .X(_05400_));
 sky130_fd_sc_hd__buf_1 _10947_ (.A(_05372_),
    .X(_05401_));
 sky130_fd_sc_hd__mux2_2 _10948_ (.A0(_05400_),
    .A1(net634),
    .S(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__buf_1 _10949_ (.A(_05402_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_2 _10950_ (.A0(_05300_),
    .A1(\rvsingle.dp.rf.rf[18][22] ),
    .S(_05401_),
    .X(_05403_));
 sky130_fd_sc_hd__buf_1 _10951_ (.A(_05403_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_2 _10952_ (.A0(_05352_),
    .A1(net271),
    .S(_05401_),
    .X(_05404_));
 sky130_fd_sc_hd__buf_1 _10953_ (.A(_05404_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_2 _10954_ (.A0(_05354_),
    .A1(net781),
    .S(_05401_),
    .X(_05405_));
 sky130_fd_sc_hd__buf_1 _10955_ (.A(_05405_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_2 _10956_ (.A0(_05304_),
    .A1(net510),
    .S(_05401_),
    .X(_05406_));
 sky130_fd_sc_hd__buf_1 _10957_ (.A(_05406_),
    .X(_00198_));
 sky130_fd_sc_hd__buf_1 _10958_ (.A(_04875_),
    .X(_05407_));
 sky130_fd_sc_hd__mux2_2 _10959_ (.A0(_05407_),
    .A1(net746),
    .S(_05401_),
    .X(_05408_));
 sky130_fd_sc_hd__buf_1 _10960_ (.A(_05408_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_2 _10961_ (.A0(_05307_),
    .A1(net594),
    .S(_05401_),
    .X(_05409_));
 sky130_fd_sc_hd__buf_1 _10962_ (.A(_05409_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_2 _10963_ (.A0(_05359_),
    .A1(net340),
    .S(_05401_),
    .X(_05410_));
 sky130_fd_sc_hd__buf_1 _10964_ (.A(_05410_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_2 _10965_ (.A0(_05266_),
    .A1(net364),
    .S(_05401_),
    .X(_05411_));
 sky130_fd_sc_hd__buf_1 _10966_ (.A(_05411_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_2 _10967_ (.A0(_05187_),
    .A1(net385),
    .S(_05401_),
    .X(_05412_));
 sky130_fd_sc_hd__buf_1 _10968_ (.A(_05412_),
    .X(_00203_));
 sky130_fd_sc_hd__inv_2 _10969_ (.A(net56),
    .Y(_05413_));
 sky130_fd_sc_hd__o21ai_2 _10970_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05368_),
    .Y(_05414_));
 sky130_fd_sc_hd__o21ai_2 _10971_ (.A1(_05413_),
    .A2(_05368_),
    .B1(_05414_),
    .Y(_00204_));
 sky130_fd_sc_hd__and3_2 _10972_ (.A(_04967_),
    .B(_04968_),
    .C(_04925_),
    .X(_05415_));
 sky130_fd_sc_hd__nor2_2 _10973_ (.A(net112),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__a21oi_2 _10974_ (.A1(_05314_),
    .A2(_05415_),
    .B1(_05416_),
    .Y(_00205_));
 sky130_fd_sc_hd__buf_1 _10975_ (.A(_04975_),
    .X(_05417_));
 sky130_fd_sc_hd__or3_2 _10976_ (.A(_04927_),
    .B(_04928_),
    .C(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__buf_1 _10977_ (.A(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__mux2_2 _10978_ (.A0(_05318_),
    .A1(\rvsingle.dp.rf.rf[31][1] ),
    .S(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__buf_1 _10979_ (.A(_05420_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_2 _10980_ (.A0(_05322_),
    .A1(net689),
    .S(_05419_),
    .X(_05421_));
 sky130_fd_sc_hd__buf_1 _10981_ (.A(_05421_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_2 _10982_ (.A0(_04755_),
    .A1(\rvsingle.dp.rf.rf[31][3] ),
    .S(_05419_),
    .X(_05422_));
 sky130_fd_sc_hd__buf_1 _10983_ (.A(_05422_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_2 _10984_ (.A0(_05377_),
    .A1(\rvsingle.dp.rf.rf[31][4] ),
    .S(_05419_),
    .X(_05423_));
 sky130_fd_sc_hd__buf_1 _10985_ (.A(_05423_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_2 _10986_ (.A0(_04765_),
    .A1(\rvsingle.dp.rf.rf[31][5] ),
    .S(_05419_),
    .X(_05424_));
 sky130_fd_sc_hd__buf_1 _10987_ (.A(_05424_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_2 _10988_ (.A0(_04770_),
    .A1(net709),
    .S(_05419_),
    .X(_05425_));
 sky130_fd_sc_hd__buf_1 _10989_ (.A(_05425_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_2 _10990_ (.A0(_05381_),
    .A1(net355),
    .S(_05419_),
    .X(_05426_));
 sky130_fd_sc_hd__buf_1 _10991_ (.A(_05426_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_2 _10992_ (.A0(_05330_),
    .A1(net737),
    .S(_05419_),
    .X(_05427_));
 sky130_fd_sc_hd__buf_1 _10993_ (.A(_05427_),
    .X(_00213_));
 sky130_fd_sc_hd__buf_1 _10994_ (.A(_04781_),
    .X(_05428_));
 sky130_fd_sc_hd__mux2_2 _10995_ (.A0(_05428_),
    .A1(net644),
    .S(_05419_),
    .X(_05429_));
 sky130_fd_sc_hd__buf_1 _10996_ (.A(_05429_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_2 _10997_ (.A0(_05385_),
    .A1(net455),
    .S(_05419_),
    .X(_05430_));
 sky130_fd_sc_hd__buf_1 _10998_ (.A(_05430_),
    .X(_00215_));
 sky130_fd_sc_hd__buf_1 _10999_ (.A(_05418_),
    .X(_05431_));
 sky130_fd_sc_hd__mux2_2 _11000_ (.A0(_05334_),
    .A1(net815),
    .S(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__buf_1 _11001_ (.A(_05432_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_2 _11002_ (.A0(_05207_),
    .A1(\rvsingle.dp.rf.rf[31][12] ),
    .S(_05431_),
    .X(_05433_));
 sky130_fd_sc_hd__buf_1 _11003_ (.A(_05433_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_2 _11004_ (.A0(_05209_),
    .A1(\rvsingle.dp.rf.rf[31][13] ),
    .S(_05431_),
    .X(_05434_));
 sky130_fd_sc_hd__buf_1 _11005_ (.A(_05434_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_2 _11006_ (.A0(_05391_),
    .A1(\rvsingle.dp.rf.rf[31][14] ),
    .S(_05431_),
    .X(_05435_));
 sky130_fd_sc_hd__buf_1 _11007_ (.A(_05435_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_2 _11008_ (.A0(_05212_),
    .A1(net812),
    .S(_05431_),
    .X(_05436_));
 sky130_fd_sc_hd__buf_1 _11009_ (.A(_05436_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_2 _11010_ (.A0(_05291_),
    .A1(\rvsingle.dp.rf.rf[31][16] ),
    .S(_05431_),
    .X(_05437_));
 sky130_fd_sc_hd__buf_1 _11011_ (.A(_05437_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_2 _11012_ (.A0(_04824_),
    .A1(\rvsingle.dp.rf.rf[31][17] ),
    .S(_05431_),
    .X(_05438_));
 sky130_fd_sc_hd__buf_1 _11013_ (.A(_05438_),
    .X(_00222_));
 sky130_fd_sc_hd__buf_1 _11014_ (.A(_04827_),
    .X(_05439_));
 sky130_fd_sc_hd__mux2_2 _11015_ (.A0(_05439_),
    .A1(\rvsingle.dp.rf.rf[31][18] ),
    .S(_05431_),
    .X(_05440_));
 sky130_fd_sc_hd__buf_1 _11016_ (.A(_05440_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_2 _11017_ (.A0(_05295_),
    .A1(\rvsingle.dp.rf.rf[31][19] ),
    .S(_05431_),
    .X(_05441_));
 sky130_fd_sc_hd__buf_1 _11018_ (.A(_05441_),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_2 _11019_ (.A0(_05398_),
    .A1(\rvsingle.dp.rf.rf[31][20] ),
    .S(_05431_),
    .X(_05442_));
 sky130_fd_sc_hd__buf_1 _11020_ (.A(_05442_),
    .X(_00225_));
 sky130_fd_sc_hd__buf_1 _11021_ (.A(_05418_),
    .X(_05443_));
 sky130_fd_sc_hd__mux2_2 _11022_ (.A0(_05400_),
    .A1(\rvsingle.dp.rf.rf[31][21] ),
    .S(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__buf_1 _11023_ (.A(_05444_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_2 _11024_ (.A0(_05300_),
    .A1(\rvsingle.dp.rf.rf[31][22] ),
    .S(_05443_),
    .X(_05445_));
 sky130_fd_sc_hd__buf_1 _11025_ (.A(_05445_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_2 _11026_ (.A0(_05352_),
    .A1(\rvsingle.dp.rf.rf[31][23] ),
    .S(_05443_),
    .X(_05446_));
 sky130_fd_sc_hd__buf_1 _11027_ (.A(_05446_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_2 _11028_ (.A0(_05354_),
    .A1(net772),
    .S(_05443_),
    .X(_05447_));
 sky130_fd_sc_hd__buf_1 _11029_ (.A(_05447_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_2 _11030_ (.A0(_05304_),
    .A1(net637),
    .S(_05443_),
    .X(_05448_));
 sky130_fd_sc_hd__buf_1 _11031_ (.A(_05448_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_2 _11032_ (.A0(_05407_),
    .A1(net502),
    .S(_05443_),
    .X(_05449_));
 sky130_fd_sc_hd__buf_1 _11033_ (.A(_05449_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_2 _11034_ (.A0(_05307_),
    .A1(net657),
    .S(_05443_),
    .X(_05450_));
 sky130_fd_sc_hd__buf_1 _11035_ (.A(_05450_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_2 _11036_ (.A0(_05359_),
    .A1(net698),
    .S(_05443_),
    .X(_05451_));
 sky130_fd_sc_hd__buf_1 _11037_ (.A(_05451_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_2 _11038_ (.A0(_05266_),
    .A1(net443),
    .S(_05443_),
    .X(_05452_));
 sky130_fd_sc_hd__buf_1 _11039_ (.A(_05452_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_2 _11040_ (.A0(_05187_),
    .A1(net426),
    .S(_05443_),
    .X(_05453_));
 sky130_fd_sc_hd__buf_1 _11041_ (.A(_05453_),
    .X(_00235_));
 sky130_fd_sc_hd__inv_2 _11042_ (.A(net81),
    .Y(_05454_));
 sky130_fd_sc_hd__o21ai_2 _11043_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05415_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21ai_2 _11044_ (.A1(_05454_),
    .A2(_05415_),
    .B1(_05455_),
    .Y(_00236_));
 sky130_fd_sc_hd__and3_2 _11045_ (.A(_04721_),
    .B(_05058_),
    .C(_05367_),
    .X(_05456_));
 sky130_fd_sc_hd__buf_1 _11046_ (.A(_05367_),
    .X(_05457_));
 sky130_fd_sc_hd__a21oi_2 _11047_ (.A1(_05145_),
    .A2(_05457_),
    .B1(net108),
    .Y(_05458_));
 sky130_fd_sc_hd__a21oi_2 _11048_ (.A1(_05314_),
    .A2(_05456_),
    .B1(_05458_),
    .Y(_00237_));
 sky130_fd_sc_hd__or4b_2 _11049_ (.A(_04919_),
    .B(_04733_),
    .C(_05371_),
    .D_N(_04737_),
    .X(_05459_));
 sky130_fd_sc_hd__buf_1 _11050_ (.A(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__mux2_2 _11051_ (.A0(_05318_),
    .A1(net471),
    .S(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__buf_1 _11052_ (.A(_05461_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_2 _11053_ (.A0(_05322_),
    .A1(net654),
    .S(_05460_),
    .X(_05462_));
 sky130_fd_sc_hd__buf_1 _11054_ (.A(_05462_),
    .X(_00239_));
 sky130_fd_sc_hd__buf_1 _11055_ (.A(_05460_),
    .X(_05463_));
 sky130_fd_sc_hd__buf_1 _11056_ (.A(_05457_),
    .X(_05464_));
 sky130_fd_sc_hd__a22o_2 _11057_ (.A1(_05463_),
    .A2(net121),
    .B1(_05156_),
    .B2(_05464_),
    .X(_00240_));
 sky130_fd_sc_hd__o311a_2 _11058_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_05061_),
    .C1(_04759_),
    .X(_05465_));
 sky130_fd_sc_hd__a22o_2 _11059_ (.A1(net198),
    .A2(_05460_),
    .B1(_05465_),
    .B2(_05464_),
    .X(_00241_));
 sky130_fd_sc_hd__a22o_2 _11060_ (.A1(_05463_),
    .A2(net159),
    .B1(_05159_),
    .B2(_05464_),
    .X(_00242_));
 sky130_fd_sc_hd__o311a_2 _11061_ (.A1(_05113_),
    .A2(_05114_),
    .A3(_05115_),
    .B1(_05061_),
    .C1(_04769_),
    .X(_05466_));
 sky130_fd_sc_hd__a22o_2 _11062_ (.A1(net54),
    .A2(_05460_),
    .B1(_05466_),
    .B2(_05464_),
    .X(_00243_));
 sky130_fd_sc_hd__a22o_2 _11063_ (.A1(_05463_),
    .A2(net135),
    .B1(_05161_),
    .B2(_05464_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_2 _11064_ (.A0(_05330_),
    .A1(net374),
    .S(_05460_),
    .X(_05467_));
 sky130_fd_sc_hd__buf_1 _11065_ (.A(_05467_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_2 _11066_ (.A0(_05428_),
    .A1(net448),
    .S(_05460_),
    .X(_05468_));
 sky130_fd_sc_hd__buf_1 _11067_ (.A(_05468_),
    .X(_00246_));
 sky130_fd_sc_hd__a22o_2 _11068_ (.A1(_05463_),
    .A2(net167),
    .B1(_05164_),
    .B2(_05464_),
    .X(_00247_));
 sky130_fd_sc_hd__buf_1 _11069_ (.A(_05459_),
    .X(_05469_));
 sky130_fd_sc_hd__mux2_2 _11070_ (.A0(_05334_),
    .A1(net595),
    .S(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__buf_1 _11071_ (.A(_05470_),
    .X(_00248_));
 sky130_fd_sc_hd__buf_1 _11072_ (.A(_05371_),
    .X(_05471_));
 sky130_fd_sc_hd__nand2_2 _11073_ (.A(_04796_),
    .B(_05145_),
    .Y(_05472_));
 sky130_fd_sc_hd__a2bb2o_2 _11074_ (.A1_N(_05471_),
    .A2_N(_05472_),
    .B1(_05463_),
    .B2(net122),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_2 _11075_ (.A0(_05209_),
    .A1(net692),
    .S(_05469_),
    .X(_05473_));
 sky130_fd_sc_hd__buf_1 _11076_ (.A(_05473_),
    .X(_00250_));
 sky130_fd_sc_hd__a2bb2o_2 _11077_ (.A1_N(_05169_),
    .A2_N(_05471_),
    .B1(_05463_),
    .B2(net158),
    .X(_00251_));
 sky130_fd_sc_hd__nand2_2 _11078_ (.A(_04814_),
    .B(_05145_),
    .Y(_05474_));
 sky130_fd_sc_hd__a2bb2o_2 _11079_ (.A1_N(_05471_),
    .A2_N(_05474_),
    .B1(_05463_),
    .B2(net183),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_2 _11080_ (.A0(_05291_),
    .A1(\rvsingle.dp.rf.rf[17][16] ),
    .S(_05469_),
    .X(_05475_));
 sky130_fd_sc_hd__buf_1 _11081_ (.A(_05475_),
    .X(_00253_));
 sky130_fd_sc_hd__buf_1 _11082_ (.A(_04823_),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_2 _11083_ (.A0(_05476_),
    .A1(net290),
    .S(_05469_),
    .X(_05477_));
 sky130_fd_sc_hd__buf_1 _11084_ (.A(_05477_),
    .X(_00254_));
 sky130_fd_sc_hd__a22o_2 _11085_ (.A1(_05463_),
    .A2(net188),
    .B1(_05174_),
    .B2(_05464_),
    .X(_00255_));
 sky130_fd_sc_hd__a2bb2o_2 _11086_ (.A1_N(_05175_),
    .A2_N(_05471_),
    .B1(_05463_),
    .B2(net137),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_2 _11087_ (.A0(_05398_),
    .A1(\rvsingle.dp.rf.rf[17][20] ),
    .S(_05469_),
    .X(_05478_));
 sky130_fd_sc_hd__buf_1 _11088_ (.A(_05478_),
    .X(_00257_));
 sky130_fd_sc_hd__a2bb2o_2 _11089_ (.A1_N(_05177_),
    .A2_N(_05471_),
    .B1(_05463_),
    .B2(net208),
    .X(_00258_));
 sky130_fd_sc_hd__a22o_2 _11090_ (.A1(_05460_),
    .A2(net162),
    .B1(_05178_),
    .B2(_05464_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_2 _11091_ (.A0(_05352_),
    .A1(\rvsingle.dp.rf.rf[17][23] ),
    .S(_05469_),
    .X(_05479_));
 sky130_fd_sc_hd__buf_1 _11092_ (.A(_05479_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_2 _11093_ (.A0(_05354_),
    .A1(\rvsingle.dp.rf.rf[17][24] ),
    .S(_05469_),
    .X(_05480_));
 sky130_fd_sc_hd__buf_1 _11094_ (.A(_05480_),
    .X(_00261_));
 sky130_fd_sc_hd__a22o_2 _11095_ (.A1(_05460_),
    .A2(net191),
    .B1(_05181_),
    .B2(_05464_),
    .X(_00262_));
 sky130_fd_sc_hd__a22o_2 _11096_ (.A1(_05460_),
    .A2(net179),
    .B1(_05182_),
    .B2(_05464_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_2 _11097_ (.A0(_05307_),
    .A1(net606),
    .S(_05469_),
    .X(_05481_));
 sky130_fd_sc_hd__buf_1 _11098_ (.A(_05481_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_2 _11099_ (.A0(_05359_),
    .A1(net408),
    .S(_05469_),
    .X(_05482_));
 sky130_fd_sc_hd__buf_1 _11100_ (.A(_05482_),
    .X(_00265_));
 sky130_fd_sc_hd__o21a_2 _11101_ (.A1(_05084_),
    .A2(_05371_),
    .B1(net652),
    .X(_05483_));
 sky130_fd_sc_hd__a31o_2 _11102_ (.A1(_04898_),
    .A2(_05183_),
    .A3(_05457_),
    .B1(_05483_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_2 _11103_ (.A0(_05187_),
    .A1(net311),
    .S(_05469_),
    .X(_05484_));
 sky130_fd_sc_hd__buf_1 _11104_ (.A(_05484_),
    .X(_00267_));
 sky130_fd_sc_hd__inv_2 _11105_ (.A(net57),
    .Y(_05485_));
 sky130_fd_sc_hd__o21ai_2 _11106_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05456_),
    .Y(_05486_));
 sky130_fd_sc_hd__o21ai_2 _11107_ (.A1(_05485_),
    .A2(_05456_),
    .B1(_05486_),
    .Y(_00268_));
 sky130_fd_sc_hd__and3_2 _11108_ (.A(_04721_),
    .B(_04924_),
    .C(_05367_),
    .X(_05487_));
 sky130_fd_sc_hd__a21oi_2 _11109_ (.A1(_05099_),
    .A2(_05457_),
    .B1(net110),
    .Y(_05488_));
 sky130_fd_sc_hd__a21oi_2 _11110_ (.A1(_05314_),
    .A2(_05487_),
    .B1(_05488_),
    .Y(_00269_));
 sky130_fd_sc_hd__or4_2 _11111_ (.A(_04737_),
    .B(_04919_),
    .C(_04733_),
    .D(_05371_),
    .X(_05489_));
 sky130_fd_sc_hd__buf_1 _11112_ (.A(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__mux2_2 _11113_ (.A0(_05318_),
    .A1(net795),
    .S(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__buf_1 _11114_ (.A(_05491_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_2 _11115_ (.A0(_05322_),
    .A1(net572),
    .S(_05490_),
    .X(_05492_));
 sky130_fd_sc_hd__buf_1 _11116_ (.A(_05492_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_2 _11117_ (.A0(_04755_),
    .A1(net702),
    .S(_05490_),
    .X(_05493_));
 sky130_fd_sc_hd__buf_1 _11118_ (.A(_05493_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_2 _11119_ (.A0(_05377_),
    .A1(net633),
    .S(_05490_),
    .X(_05494_));
 sky130_fd_sc_hd__buf_1 _11120_ (.A(_05494_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_2 _11121_ (.A0(_04765_),
    .A1(\rvsingle.dp.rf.rf[16][5] ),
    .S(_05490_),
    .X(_05495_));
 sky130_fd_sc_hd__buf_1 _11122_ (.A(_05495_),
    .X(_00274_));
 sky130_fd_sc_hd__buf_1 _11123_ (.A(_04769_),
    .X(_05496_));
 sky130_fd_sc_hd__mux2_2 _11124_ (.A0(_05496_),
    .A1(\rvsingle.dp.rf.rf[16][6] ),
    .S(_05490_),
    .X(_05497_));
 sky130_fd_sc_hd__buf_1 _11125_ (.A(_05497_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_2 _11126_ (.A0(_05381_),
    .A1(net399),
    .S(_05490_),
    .X(_05498_));
 sky130_fd_sc_hd__buf_1 _11127_ (.A(_05498_),
    .X(_00276_));
 sky130_fd_sc_hd__buf_1 _11128_ (.A(_05489_),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_2 _11129_ (.A0(_05330_),
    .A1(\rvsingle.dp.rf.rf[16][8] ),
    .S(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__buf_1 _11130_ (.A(_05500_),
    .X(_00277_));
 sky130_fd_sc_hd__buf_1 _11131_ (.A(_05367_),
    .X(_05501_));
 sky130_fd_sc_hd__a22o_2 _11132_ (.A1(_05490_),
    .A2(net123),
    .B1(_05116_),
    .B2(_05501_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_2 _11133_ (.A0(_05385_),
    .A1(net533),
    .S(_05499_),
    .X(_05502_));
 sky130_fd_sc_hd__buf_1 _11134_ (.A(_05502_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_2 _11135_ (.A0(_05334_),
    .A1(net432),
    .S(_05499_),
    .X(_05503_));
 sky130_fd_sc_hd__buf_1 _11136_ (.A(_05503_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_2 _11137_ (.A0(_05207_),
    .A1(\rvsingle.dp.rf.rf[16][12] ),
    .S(_05499_),
    .X(_05504_));
 sky130_fd_sc_hd__buf_1 _11138_ (.A(_05504_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_2 _11139_ (.A0(_05209_),
    .A1(\rvsingle.dp.rf.rf[16][13] ),
    .S(_05499_),
    .X(_05505_));
 sky130_fd_sc_hd__buf_1 _11140_ (.A(_05505_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_2 _11141_ (.A0(_05391_),
    .A1(\rvsingle.dp.rf.rf[16][14] ),
    .S(_05499_),
    .X(_05506_));
 sky130_fd_sc_hd__buf_1 _11142_ (.A(_05506_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_2 _11143_ (.A0(_05212_),
    .A1(\rvsingle.dp.rf.rf[16][15] ),
    .S(_05499_),
    .X(_05507_));
 sky130_fd_sc_hd__buf_1 _11144_ (.A(_05507_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_2 _11145_ (.A0(_05291_),
    .A1(net522),
    .S(_05499_),
    .X(_05508_));
 sky130_fd_sc_hd__buf_1 _11146_ (.A(_05508_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_2 _11147_ (.A0(_05476_),
    .A1(net658),
    .S(_05499_),
    .X(_05509_));
 sky130_fd_sc_hd__buf_1 _11148_ (.A(_05509_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_2 _11149_ (.A0(_05439_),
    .A1(\rvsingle.dp.rf.rf[16][18] ),
    .S(_05499_),
    .X(_05510_));
 sky130_fd_sc_hd__buf_1 _11150_ (.A(_05510_),
    .X(_00287_));
 sky130_fd_sc_hd__buf_1 _11151_ (.A(_05489_),
    .X(_05511_));
 sky130_fd_sc_hd__mux2_2 _11152_ (.A0(_05295_),
    .A1(net673),
    .S(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__buf_1 _11153_ (.A(_05512_),
    .X(_00288_));
 sky130_fd_sc_hd__or4b_2 _11154_ (.A(_04967_),
    .B(_04968_),
    .C(_04976_),
    .D_N(_04839_),
    .X(_05513_));
 sky130_fd_sc_hd__o2bb2ai_2 _11155_ (.A1_N(_05490_),
    .A2_N(net16),
    .B1(_05371_),
    .B2(_05513_),
    .Y(_00289_));
 sky130_fd_sc_hd__mux2_2 _11156_ (.A0(_05400_),
    .A1(net793),
    .S(_05511_),
    .X(_05514_));
 sky130_fd_sc_hd__buf_1 _11157_ (.A(_05514_),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_2 _11158_ (.A0(_05300_),
    .A1(net220),
    .S(_05511_),
    .X(_05515_));
 sky130_fd_sc_hd__buf_1 _11159_ (.A(_05515_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_2 _11160_ (.A0(_05352_),
    .A1(net460),
    .S(_05511_),
    .X(_05516_));
 sky130_fd_sc_hd__buf_1 _11161_ (.A(_05516_),
    .X(_00292_));
 sky130_fd_sc_hd__a22o_2 _11162_ (.A1(_05490_),
    .A2(net197),
    .B1(_05133_),
    .B2(_05501_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_2 _11163_ (.A0(_05304_),
    .A1(net335),
    .S(_05511_),
    .X(_05517_));
 sky130_fd_sc_hd__buf_1 _11164_ (.A(_05517_),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_2 _11165_ (.A0(_05407_),
    .A1(\rvsingle.dp.rf.rf[16][26] ),
    .S(_05511_),
    .X(_05518_));
 sky130_fd_sc_hd__buf_1 _11166_ (.A(_05518_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_2 _11167_ (.A0(_05307_),
    .A1(net451),
    .S(_05511_),
    .X(_05519_));
 sky130_fd_sc_hd__buf_1 _11168_ (.A(_05519_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_2 _11169_ (.A0(_05359_),
    .A1(net351),
    .S(_05511_),
    .X(_05520_));
 sky130_fd_sc_hd__buf_1 _11170_ (.A(_05520_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_2 _11171_ (.A0(_05266_),
    .A1(net429),
    .S(_05511_),
    .X(_05521_));
 sky130_fd_sc_hd__buf_1 _11172_ (.A(_05521_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_2 _11173_ (.A0(_05187_),
    .A1(net361),
    .S(_05511_),
    .X(_05522_));
 sky130_fd_sc_hd__buf_1 _11174_ (.A(_05522_),
    .X(_00299_));
 sky130_fd_sc_hd__inv_2 _11175_ (.A(net46),
    .Y(_05523_));
 sky130_fd_sc_hd__o21ai_2 _11176_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05487_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21ai_2 _11177_ (.A1(_05523_),
    .A2(_05487_),
    .B1(_05524_),
    .Y(_00300_));
 sky130_fd_sc_hd__and4_2 _11178_ (.A(_04916_),
    .B(_04918_),
    .C(_04922_),
    .D(_05058_),
    .X(_05525_));
 sky130_fd_sc_hd__a21oi_2 _11179_ (.A1(_04925_),
    .A2(_05061_),
    .B1(net74),
    .Y(_05526_));
 sky130_fd_sc_hd__a21oi_2 _11180_ (.A1(_05314_),
    .A2(_05525_),
    .B1(_05526_),
    .Y(_00301_));
 sky130_fd_sc_hd__or4b_2 _11181_ (.A(_04919_),
    .B(_04927_),
    .C(_04928_),
    .D_N(_04738_),
    .X(_05527_));
 sky130_fd_sc_hd__buf_1 _11182_ (.A(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_2 _11183_ (.A0(_05318_),
    .A1(net766),
    .S(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__buf_1 _11184_ (.A(_05529_),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_2 _11185_ (.A0(_05322_),
    .A1(net805),
    .S(_05528_),
    .X(_05530_));
 sky130_fd_sc_hd__buf_1 _11186_ (.A(_05530_),
    .X(_00303_));
 sky130_fd_sc_hd__buf_1 _11187_ (.A(_04754_),
    .X(_05531_));
 sky130_fd_sc_hd__mux2_2 _11188_ (.A0(_05531_),
    .A1(net816),
    .S(_05528_),
    .X(_05532_));
 sky130_fd_sc_hd__buf_1 _11189_ (.A(_05532_),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_2 _11190_ (.A0(_05377_),
    .A1(net740),
    .S(_05528_),
    .X(_05533_));
 sky130_fd_sc_hd__buf_1 _11191_ (.A(_05533_),
    .X(_00305_));
 sky130_fd_sc_hd__buf_1 _11192_ (.A(_04764_),
    .X(_05534_));
 sky130_fd_sc_hd__mux2_2 _11193_ (.A0(_05534_),
    .A1(net752),
    .S(_05528_),
    .X(_05535_));
 sky130_fd_sc_hd__buf_1 _11194_ (.A(_05535_),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_2 _11195_ (.A0(_05496_),
    .A1(net757),
    .S(_05528_),
    .X(_05536_));
 sky130_fd_sc_hd__buf_1 _11196_ (.A(_05536_),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_2 _11197_ (.A0(_05381_),
    .A1(net444),
    .S(_05528_),
    .X(_05537_));
 sky130_fd_sc_hd__buf_1 _11198_ (.A(_05537_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_2 _11199_ (.A0(_05330_),
    .A1(net419),
    .S(_05528_),
    .X(_05538_));
 sky130_fd_sc_hd__buf_1 _11200_ (.A(_05538_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_2 _11201_ (.A0(_05428_),
    .A1(net404),
    .S(_05528_),
    .X(_05539_));
 sky130_fd_sc_hd__buf_1 _11202_ (.A(_05539_),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_2 _11203_ (.A0(_05385_),
    .A1(net431),
    .S(_05528_),
    .X(_05540_));
 sky130_fd_sc_hd__buf_1 _11204_ (.A(_05540_),
    .X(_00311_));
 sky130_fd_sc_hd__buf_1 _11205_ (.A(_05527_),
    .X(_05541_));
 sky130_fd_sc_hd__mux2_2 _11206_ (.A0(_05334_),
    .A1(net796),
    .S(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__buf_1 _11207_ (.A(_05542_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_2 _11208_ (.A0(_05207_),
    .A1(net534),
    .S(_05541_),
    .X(_05543_));
 sky130_fd_sc_hd__buf_1 _11209_ (.A(_05543_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_2 _11210_ (.A0(_05209_),
    .A1(\rvsingle.dp.rf.rf[29][13] ),
    .S(_05541_),
    .X(_05544_));
 sky130_fd_sc_hd__buf_1 _11211_ (.A(_05544_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_2 _11212_ (.A0(_05391_),
    .A1(\rvsingle.dp.rf.rf[29][14] ),
    .S(_05541_),
    .X(_05545_));
 sky130_fd_sc_hd__buf_1 _11213_ (.A(_05545_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_2 _11214_ (.A0(_05212_),
    .A1(\rvsingle.dp.rf.rf[29][15] ),
    .S(_05541_),
    .X(_05546_));
 sky130_fd_sc_hd__buf_1 _11215_ (.A(_05546_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_2 _11216_ (.A0(_05291_),
    .A1(\rvsingle.dp.rf.rf[29][16] ),
    .S(_05541_),
    .X(_05547_));
 sky130_fd_sc_hd__buf_1 _11217_ (.A(_05547_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_2 _11218_ (.A0(_05476_),
    .A1(net668),
    .S(_05541_),
    .X(_05548_));
 sky130_fd_sc_hd__buf_1 _11219_ (.A(_05548_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_2 _11220_ (.A0(_05439_),
    .A1(\rvsingle.dp.rf.rf[29][18] ),
    .S(_05541_),
    .X(_05549_));
 sky130_fd_sc_hd__buf_1 _11221_ (.A(_05549_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_2 _11222_ (.A0(_05295_),
    .A1(\rvsingle.dp.rf.rf[29][19] ),
    .S(_05541_),
    .X(_05550_));
 sky130_fd_sc_hd__buf_1 _11223_ (.A(_05550_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_2 _11224_ (.A0(_05398_),
    .A1(net705),
    .S(_05541_),
    .X(_05551_));
 sky130_fd_sc_hd__buf_1 _11225_ (.A(_05551_),
    .X(_00321_));
 sky130_fd_sc_hd__buf_1 _11226_ (.A(_05527_),
    .X(_05552_));
 sky130_fd_sc_hd__mux2_2 _11227_ (.A0(_05400_),
    .A1(\rvsingle.dp.rf.rf[29][21] ),
    .S(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__buf_1 _11228_ (.A(_05553_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_2 _11229_ (.A0(_05300_),
    .A1(\rvsingle.dp.rf.rf[29][22] ),
    .S(_05552_),
    .X(_05554_));
 sky130_fd_sc_hd__buf_1 _11230_ (.A(_05554_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_2 _11231_ (.A0(_05352_),
    .A1(\rvsingle.dp.rf.rf[29][23] ),
    .S(_05552_),
    .X(_05555_));
 sky130_fd_sc_hd__buf_1 _11232_ (.A(_05555_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_2 _11233_ (.A0(_05354_),
    .A1(\rvsingle.dp.rf.rf[29][24] ),
    .S(_05552_),
    .X(_05556_));
 sky130_fd_sc_hd__buf_1 _11234_ (.A(_05556_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_2 _11235_ (.A0(_05304_),
    .A1(net800),
    .S(_05552_),
    .X(_05557_));
 sky130_fd_sc_hd__buf_1 _11236_ (.A(_05557_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_2 _11237_ (.A0(_05407_),
    .A1(net603),
    .S(_05552_),
    .X(_05558_));
 sky130_fd_sc_hd__buf_1 _11238_ (.A(_05558_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_2 _11239_ (.A0(_05307_),
    .A1(net621),
    .S(_05552_),
    .X(_05559_));
 sky130_fd_sc_hd__buf_1 _11240_ (.A(_05559_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_2 _11241_ (.A0(_05359_),
    .A1(net291),
    .S(_05552_),
    .X(_05560_));
 sky130_fd_sc_hd__buf_1 _11242_ (.A(_05560_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_2 _11243_ (.A0(_05266_),
    .A1(net328),
    .S(_05552_),
    .X(_05561_));
 sky130_fd_sc_hd__buf_1 _11244_ (.A(_05561_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_2 _11245_ (.A0(_05187_),
    .A1(net302),
    .S(_05552_),
    .X(_05562_));
 sky130_fd_sc_hd__buf_1 _11246_ (.A(_05562_),
    .X(_00331_));
 sky130_fd_sc_hd__inv_2 _11247_ (.A(net80),
    .Y(_05563_));
 sky130_fd_sc_hd__o21ai_2 _11248_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05525_),
    .Y(_05564_));
 sky130_fd_sc_hd__o21ai_2 _11249_ (.A1(_05563_),
    .A2(_05525_),
    .B1(_05564_),
    .Y(_00332_));
 sky130_fd_sc_hd__or3b_2 _11250_ (.A(_04928_),
    .B(_04722_),
    .C_N(_04723_),
    .X(_05565_));
 sky130_fd_sc_hd__nor2_2 _11251_ (.A(_05417_),
    .B(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__nor2_2 _11252_ (.A(net142),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__a21oi_2 _11253_ (.A1(_05314_),
    .A2(_05566_),
    .B1(_05567_),
    .Y(_00333_));
 sky130_fd_sc_hd__or2_2 _11254_ (.A(_05417_),
    .B(_05565_),
    .X(_05568_));
 sky130_fd_sc_hd__buf_1 _11255_ (.A(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__mux2_2 _11256_ (.A0(_05318_),
    .A1(\rvsingle.dp.rf.rf[15][1] ),
    .S(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__buf_1 _11257_ (.A(_05570_),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_2 _11258_ (.A0(_05322_),
    .A1(\rvsingle.dp.rf.rf[15][2] ),
    .S(_05569_),
    .X(_05571_));
 sky130_fd_sc_hd__buf_1 _11259_ (.A(_05571_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_2 _11260_ (.A0(_05531_),
    .A1(\rvsingle.dp.rf.rf[15][3] ),
    .S(_05569_),
    .X(_05572_));
 sky130_fd_sc_hd__buf_1 _11261_ (.A(_05572_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_2 _11262_ (.A0(_05377_),
    .A1(\rvsingle.dp.rf.rf[15][4] ),
    .S(_05569_),
    .X(_05573_));
 sky130_fd_sc_hd__buf_1 _11263_ (.A(_05573_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_2 _11264_ (.A0(_05534_),
    .A1(net741),
    .S(_05569_),
    .X(_05574_));
 sky130_fd_sc_hd__buf_1 _11265_ (.A(_05574_),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_2 _11266_ (.A0(_05496_),
    .A1(net646),
    .S(_05569_),
    .X(_05575_));
 sky130_fd_sc_hd__buf_1 _11267_ (.A(_05575_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_2 _11268_ (.A0(_05381_),
    .A1(net724),
    .S(_05569_),
    .X(_05576_));
 sky130_fd_sc_hd__buf_1 _11269_ (.A(_05576_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_2 _11270_ (.A0(_05330_),
    .A1(net806),
    .S(_05569_),
    .X(_05577_));
 sky130_fd_sc_hd__buf_1 _11271_ (.A(_05577_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_2 _11272_ (.A0(_05428_),
    .A1(net501),
    .S(_05569_),
    .X(_05578_));
 sky130_fd_sc_hd__buf_1 _11273_ (.A(_05578_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_2 _11274_ (.A0(_05385_),
    .A1(\rvsingle.dp.rf.rf[15][10] ),
    .S(_05569_),
    .X(_05579_));
 sky130_fd_sc_hd__buf_1 _11275_ (.A(_05579_),
    .X(_00343_));
 sky130_fd_sc_hd__buf_1 _11276_ (.A(_05568_),
    .X(_05580_));
 sky130_fd_sc_hd__mux2_2 _11277_ (.A0(_05334_),
    .A1(net717),
    .S(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__buf_1 _11278_ (.A(_05581_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_2 _11279_ (.A0(_05207_),
    .A1(net438),
    .S(_05580_),
    .X(_05582_));
 sky130_fd_sc_hd__buf_1 _11280_ (.A(_05582_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_2 _11281_ (.A0(_05209_),
    .A1(\rvsingle.dp.rf.rf[15][13] ),
    .S(_05580_),
    .X(_05583_));
 sky130_fd_sc_hd__buf_1 _11282_ (.A(_05583_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_2 _11283_ (.A0(_05391_),
    .A1(\rvsingle.dp.rf.rf[15][14] ),
    .S(_05580_),
    .X(_05584_));
 sky130_fd_sc_hd__buf_1 _11284_ (.A(_05584_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_2 _11285_ (.A0(_05212_),
    .A1(net744),
    .S(_05580_),
    .X(_05585_));
 sky130_fd_sc_hd__buf_1 _11286_ (.A(_05585_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_2 _11287_ (.A0(_05291_),
    .A1(net803),
    .S(_05580_),
    .X(_05586_));
 sky130_fd_sc_hd__buf_1 _11288_ (.A(_05586_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_2 _11289_ (.A0(_05476_),
    .A1(net544),
    .S(_05580_),
    .X(_05587_));
 sky130_fd_sc_hd__buf_1 _11290_ (.A(_05587_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_2 _11291_ (.A0(_05439_),
    .A1(\rvsingle.dp.rf.rf[15][18] ),
    .S(_05580_),
    .X(_05588_));
 sky130_fd_sc_hd__buf_1 _11292_ (.A(_05588_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_2 _11293_ (.A0(_05295_),
    .A1(net729),
    .S(_05580_),
    .X(_05589_));
 sky130_fd_sc_hd__buf_1 _11294_ (.A(_05589_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_2 _11295_ (.A0(_05398_),
    .A1(net788),
    .S(_05580_),
    .X(_05590_));
 sky130_fd_sc_hd__buf_1 _11296_ (.A(_05590_),
    .X(_00353_));
 sky130_fd_sc_hd__buf_1 _11297_ (.A(_05568_),
    .X(_05591_));
 sky130_fd_sc_hd__mux2_2 _11298_ (.A0(_05400_),
    .A1(\rvsingle.dp.rf.rf[15][21] ),
    .S(_05591_),
    .X(_05592_));
 sky130_fd_sc_hd__buf_1 _11299_ (.A(_05592_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_2 _11300_ (.A0(_05300_),
    .A1(\rvsingle.dp.rf.rf[15][22] ),
    .S(_05591_),
    .X(_05593_));
 sky130_fd_sc_hd__buf_1 _11301_ (.A(_05593_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_2 _11302_ (.A0(_05352_),
    .A1(\rvsingle.dp.rf.rf[15][23] ),
    .S(_05591_),
    .X(_05594_));
 sky130_fd_sc_hd__buf_1 _11303_ (.A(_05594_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_2 _11304_ (.A0(_05354_),
    .A1(\rvsingle.dp.rf.rf[15][24] ),
    .S(_05591_),
    .X(_05595_));
 sky130_fd_sc_hd__buf_1 _11305_ (.A(_05595_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_2 _11306_ (.A0(_05304_),
    .A1(\rvsingle.dp.rf.rf[15][25] ),
    .S(_05591_),
    .X(_05596_));
 sky130_fd_sc_hd__buf_1 _11307_ (.A(_05596_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_2 _11308_ (.A0(_05407_),
    .A1(net508),
    .S(_05591_),
    .X(_05597_));
 sky130_fd_sc_hd__buf_1 _11309_ (.A(_05597_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_2 _11310_ (.A0(_05307_),
    .A1(\rvsingle.dp.rf.rf[15][27] ),
    .S(_05591_),
    .X(_05598_));
 sky130_fd_sc_hd__buf_1 _11311_ (.A(_05598_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_2 _11312_ (.A0(_05359_),
    .A1(net449),
    .S(_05591_),
    .X(_05599_));
 sky130_fd_sc_hd__buf_1 _11313_ (.A(_05599_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_2 _11314_ (.A0(_05266_),
    .A1(net440),
    .S(_05591_),
    .X(_05600_));
 sky130_fd_sc_hd__buf_1 _11315_ (.A(_05600_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_2 _11316_ (.A0(_05187_),
    .A1(net407),
    .S(_05591_),
    .X(_05601_));
 sky130_fd_sc_hd__buf_1 _11317_ (.A(_05601_),
    .X(_00363_));
 sky130_fd_sc_hd__inv_2 _11318_ (.A(net70),
    .Y(_05602_));
 sky130_fd_sc_hd__o21ai_2 _11319_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05566_),
    .Y(_05603_));
 sky130_fd_sc_hd__o21ai_2 _11320_ (.A1(_05602_),
    .A2(_05566_),
    .B1(_05603_),
    .Y(_00364_));
 sky130_fd_sc_hd__and4b_2 _11321_ (.A_N(_04916_),
    .B(_04918_),
    .C(_04728_),
    .D(_04922_),
    .X(_05604_));
 sky130_fd_sc_hd__nor2_2 _11322_ (.A(net124),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__a21oi_2 _11323_ (.A1(_05314_),
    .A2(_05604_),
    .B1(_05605_),
    .Y(_00365_));
 sky130_fd_sc_hd__or3b_2 _11324_ (.A(_05565_),
    .B(_04738_),
    .C_N(_04739_),
    .X(_05606_));
 sky130_fd_sc_hd__buf_1 _11325_ (.A(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__mux2_2 _11326_ (.A0(_05318_),
    .A1(net701),
    .S(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__buf_1 _11327_ (.A(_05608_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_2 _11328_ (.A0(_05322_),
    .A1(net473),
    .S(_05607_),
    .X(_05609_));
 sky130_fd_sc_hd__buf_1 _11329_ (.A(_05609_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_2 _11330_ (.A0(_05531_),
    .A1(\rvsingle.dp.rf.rf[14][3] ),
    .S(_05607_),
    .X(_05610_));
 sky130_fd_sc_hd__buf_1 _11331_ (.A(_05610_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_2 _11332_ (.A0(_05377_),
    .A1(net590),
    .S(_05607_),
    .X(_05611_));
 sky130_fd_sc_hd__buf_1 _11333_ (.A(_05611_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_2 _11334_ (.A0(_05534_),
    .A1(\rvsingle.dp.rf.rf[14][5] ),
    .S(_05607_),
    .X(_05612_));
 sky130_fd_sc_hd__buf_1 _11335_ (.A(_05612_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_2 _11336_ (.A0(_05496_),
    .A1(net410),
    .S(_05607_),
    .X(_05613_));
 sky130_fd_sc_hd__buf_1 _11337_ (.A(_05613_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_2 _11338_ (.A0(_05381_),
    .A1(\rvsingle.dp.rf.rf[14][7] ),
    .S(_05607_),
    .X(_05614_));
 sky130_fd_sc_hd__buf_1 _11339_ (.A(_05614_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_2 _11340_ (.A0(_05330_),
    .A1(net708),
    .S(_05607_),
    .X(_05615_));
 sky130_fd_sc_hd__buf_1 _11341_ (.A(_05615_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_2 _11342_ (.A0(_05428_),
    .A1(net495),
    .S(_05607_),
    .X(_05616_));
 sky130_fd_sc_hd__buf_1 _11343_ (.A(_05616_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_2 _11344_ (.A0(_05385_),
    .A1(\rvsingle.dp.rf.rf[14][10] ),
    .S(_05607_),
    .X(_05617_));
 sky130_fd_sc_hd__buf_1 _11345_ (.A(_05617_),
    .X(_00375_));
 sky130_fd_sc_hd__buf_1 _11346_ (.A(_05606_),
    .X(_05618_));
 sky130_fd_sc_hd__mux2_2 _11347_ (.A0(_05334_),
    .A1(net468),
    .S(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__buf_1 _11348_ (.A(_05619_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_2 _11349_ (.A0(_05207_),
    .A1(net776),
    .S(_05618_),
    .X(_05620_));
 sky130_fd_sc_hd__buf_1 _11350_ (.A(_05620_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_2 _11351_ (.A0(_05209_),
    .A1(\rvsingle.dp.rf.rf[14][13] ),
    .S(_05618_),
    .X(_05621_));
 sky130_fd_sc_hd__buf_1 _11352_ (.A(_05621_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_2 _11353_ (.A0(_05391_),
    .A1(net604),
    .S(_05618_),
    .X(_05622_));
 sky130_fd_sc_hd__buf_1 _11354_ (.A(_05622_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_2 _11355_ (.A0(_05212_),
    .A1(net761),
    .S(_05618_),
    .X(_05623_));
 sky130_fd_sc_hd__buf_1 _11356_ (.A(_05623_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_2 _11357_ (.A0(_05291_),
    .A1(\rvsingle.dp.rf.rf[14][16] ),
    .S(_05618_),
    .X(_05624_));
 sky130_fd_sc_hd__buf_1 _11358_ (.A(_05624_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_2 _11359_ (.A0(_05476_),
    .A1(net785),
    .S(_05618_),
    .X(_05625_));
 sky130_fd_sc_hd__buf_1 _11360_ (.A(_05625_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_2 _11361_ (.A0(_05439_),
    .A1(net618),
    .S(_05618_),
    .X(_05626_));
 sky130_fd_sc_hd__buf_1 _11362_ (.A(_05626_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_2 _11363_ (.A0(_05295_),
    .A1(net725),
    .S(_05618_),
    .X(_05627_));
 sky130_fd_sc_hd__buf_1 _11364_ (.A(_05627_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_2 _11365_ (.A0(_05398_),
    .A1(\rvsingle.dp.rf.rf[14][20] ),
    .S(_05618_),
    .X(_05628_));
 sky130_fd_sc_hd__buf_1 _11366_ (.A(_05628_),
    .X(_00385_));
 sky130_fd_sc_hd__buf_1 _11367_ (.A(_05606_),
    .X(_05629_));
 sky130_fd_sc_hd__mux2_2 _11368_ (.A0(_05400_),
    .A1(net810),
    .S(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__buf_1 _11369_ (.A(_05630_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_2 _11370_ (.A0(_05300_),
    .A1(\rvsingle.dp.rf.rf[14][22] ),
    .S(_05629_),
    .X(_05631_));
 sky130_fd_sc_hd__buf_1 _11371_ (.A(_05631_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_2 _11372_ (.A0(_05352_),
    .A1(\rvsingle.dp.rf.rf[14][23] ),
    .S(_05629_),
    .X(_05632_));
 sky130_fd_sc_hd__buf_1 _11373_ (.A(_05632_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_2 _11374_ (.A0(_05354_),
    .A1(\rvsingle.dp.rf.rf[14][24] ),
    .S(_05629_),
    .X(_05633_));
 sky130_fd_sc_hd__buf_1 _11375_ (.A(_05633_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_2 _11376_ (.A0(_05304_),
    .A1(net458),
    .S(_05629_),
    .X(_05634_));
 sky130_fd_sc_hd__buf_1 _11377_ (.A(_05634_),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_2 _11378_ (.A0(_05407_),
    .A1(net512),
    .S(_05629_),
    .X(_05635_));
 sky130_fd_sc_hd__buf_1 _11379_ (.A(_05635_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_2 _11380_ (.A0(_05307_),
    .A1(net728),
    .S(_05629_),
    .X(_05636_));
 sky130_fd_sc_hd__buf_1 _11381_ (.A(_05636_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_2 _11382_ (.A0(_05359_),
    .A1(net427),
    .S(_05629_),
    .X(_05637_));
 sky130_fd_sc_hd__buf_1 _11383_ (.A(_05637_),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_2 _11384_ (.A0(_05266_),
    .A1(net459),
    .S(_05629_),
    .X(_05638_));
 sky130_fd_sc_hd__buf_1 _11385_ (.A(_05638_),
    .X(_00394_));
 sky130_fd_sc_hd__buf_1 _11386_ (.A(_04903_),
    .X(_05639_));
 sky130_fd_sc_hd__mux2_2 _11387_ (.A0(_05639_),
    .A1(net295),
    .S(_05629_),
    .X(_05640_));
 sky130_fd_sc_hd__buf_1 _11388_ (.A(_05640_),
    .X(_00395_));
 sky130_fd_sc_hd__inv_2 _11389_ (.A(net71),
    .Y(_05641_));
 sky130_fd_sc_hd__o21ai_2 _11390_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05604_),
    .Y(_05642_));
 sky130_fd_sc_hd__o21ai_2 _11391_ (.A1(_05641_),
    .A2(_05604_),
    .B1(_05642_),
    .Y(_00396_));
 sky130_fd_sc_hd__and4b_2 _11392_ (.A_N(_04916_),
    .B(_04918_),
    .C(_04922_),
    .D(_05058_),
    .X(_05643_));
 sky130_fd_sc_hd__nor2_2 _11393_ (.A(net178),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__a21oi_2 _11394_ (.A1(_05314_),
    .A2(_05643_),
    .B1(_05644_),
    .Y(_00397_));
 sky130_fd_sc_hd__or3b_2 _11395_ (.A(_04739_),
    .B(_05565_),
    .C_N(_04738_),
    .X(_05645_));
 sky130_fd_sc_hd__buf_1 _11396_ (.A(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__mux2_2 _11397_ (.A0(_05318_),
    .A1(\rvsingle.dp.rf.rf[13][1] ),
    .S(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__buf_1 _11398_ (.A(_05647_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_2 _11399_ (.A0(_05322_),
    .A1(\rvsingle.dp.rf.rf[13][2] ),
    .S(_05646_),
    .X(_05648_));
 sky130_fd_sc_hd__buf_1 _11400_ (.A(_05648_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_2 _11401_ (.A0(_05531_),
    .A1(\rvsingle.dp.rf.rf[13][3] ),
    .S(_05646_),
    .X(_05649_));
 sky130_fd_sc_hd__buf_1 _11402_ (.A(_05649_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_2 _11403_ (.A0(_05377_),
    .A1(\rvsingle.dp.rf.rf[13][4] ),
    .S(_05646_),
    .X(_05650_));
 sky130_fd_sc_hd__buf_1 _11404_ (.A(_05650_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_2 _11405_ (.A0(_05534_),
    .A1(\rvsingle.dp.rf.rf[13][5] ),
    .S(_05646_),
    .X(_05651_));
 sky130_fd_sc_hd__buf_1 _11406_ (.A(_05651_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_2 _11407_ (.A0(_05496_),
    .A1(net509),
    .S(_05646_),
    .X(_05652_));
 sky130_fd_sc_hd__buf_1 _11408_ (.A(_05652_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_2 _11409_ (.A0(_05381_),
    .A1(net753),
    .S(_05646_),
    .X(_05653_));
 sky130_fd_sc_hd__buf_1 _11410_ (.A(_05653_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_2 _11411_ (.A0(_05330_),
    .A1(net726),
    .S(_05646_),
    .X(_05654_));
 sky130_fd_sc_hd__buf_1 _11412_ (.A(_05654_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_2 _11413_ (.A0(_05428_),
    .A1(net484),
    .S(_05646_),
    .X(_05655_));
 sky130_fd_sc_hd__buf_1 _11414_ (.A(_05655_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_2 _11415_ (.A0(_05385_),
    .A1(\rvsingle.dp.rf.rf[13][10] ),
    .S(_05646_),
    .X(_05656_));
 sky130_fd_sc_hd__buf_1 _11416_ (.A(_05656_),
    .X(_00407_));
 sky130_fd_sc_hd__buf_1 _11417_ (.A(_05645_),
    .X(_05657_));
 sky130_fd_sc_hd__mux2_2 _11418_ (.A0(_05334_),
    .A1(net640),
    .S(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__buf_1 _11419_ (.A(_05658_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_2 _11420_ (.A0(_05207_),
    .A1(net367),
    .S(_05657_),
    .X(_05659_));
 sky130_fd_sc_hd__buf_1 _11421_ (.A(_05659_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_2 _11422_ (.A0(_04801_),
    .A1(net488),
    .S(_05657_),
    .X(_05660_));
 sky130_fd_sc_hd__buf_1 _11423_ (.A(_05660_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_2 _11424_ (.A0(_05391_),
    .A1(net697),
    .S(_05657_),
    .X(_05661_));
 sky130_fd_sc_hd__buf_1 _11425_ (.A(_05661_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_2 _11426_ (.A0(_05212_),
    .A1(net720),
    .S(_05657_),
    .X(_05662_));
 sky130_fd_sc_hd__buf_1 _11427_ (.A(_05662_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_2 _11428_ (.A0(_05291_),
    .A1(net723),
    .S(_05657_),
    .X(_05663_));
 sky130_fd_sc_hd__buf_1 _11429_ (.A(_05663_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_2 _11430_ (.A0(_05476_),
    .A1(net611),
    .S(_05657_),
    .X(_05664_));
 sky130_fd_sc_hd__buf_1 _11431_ (.A(_05664_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_2 _11432_ (.A0(_05439_),
    .A1(net713),
    .S(_05657_),
    .X(_05665_));
 sky130_fd_sc_hd__buf_1 _11433_ (.A(_05665_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_2 _11434_ (.A0(_05295_),
    .A1(net559),
    .S(_05657_),
    .X(_05666_));
 sky130_fd_sc_hd__buf_1 _11435_ (.A(_05666_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_2 _11436_ (.A0(_05398_),
    .A1(net801),
    .S(_05657_),
    .X(_05667_));
 sky130_fd_sc_hd__buf_1 _11437_ (.A(_05667_),
    .X(_00417_));
 sky130_fd_sc_hd__buf_1 _11438_ (.A(_05645_),
    .X(_05668_));
 sky130_fd_sc_hd__mux2_2 _11439_ (.A0(_05400_),
    .A1(\rvsingle.dp.rf.rf[13][21] ),
    .S(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__buf_1 _11440_ (.A(_05669_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_2 _11441_ (.A0(_05300_),
    .A1(\rvsingle.dp.rf.rf[13][22] ),
    .S(_05668_),
    .X(_05670_));
 sky130_fd_sc_hd__buf_1 _11442_ (.A(_05670_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_2 _11443_ (.A0(_05352_),
    .A1(\rvsingle.dp.rf.rf[13][23] ),
    .S(_05668_),
    .X(_05671_));
 sky130_fd_sc_hd__buf_1 _11444_ (.A(_05671_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_2 _11445_ (.A0(_05354_),
    .A1(\rvsingle.dp.rf.rf[13][24] ),
    .S(_05668_),
    .X(_05672_));
 sky130_fd_sc_hd__buf_1 _11446_ (.A(_05672_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_2 _11447_ (.A0(_05304_),
    .A1(\rvsingle.dp.rf.rf[13][25] ),
    .S(_05668_),
    .X(_05673_));
 sky130_fd_sc_hd__buf_1 _11448_ (.A(_05673_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_2 _11449_ (.A0(_05407_),
    .A1(net645),
    .S(_05668_),
    .X(_05674_));
 sky130_fd_sc_hd__buf_1 _11450_ (.A(_05674_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_2 _11451_ (.A0(_05307_),
    .A1(\rvsingle.dp.rf.rf[13][27] ),
    .S(_05668_),
    .X(_05675_));
 sky130_fd_sc_hd__buf_1 _11452_ (.A(_05675_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_2 _11453_ (.A0(_05359_),
    .A1(net465),
    .S(_05668_),
    .X(_05676_));
 sky130_fd_sc_hd__buf_1 _11454_ (.A(_05676_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_2 _11455_ (.A0(_05266_),
    .A1(net503),
    .S(_05668_),
    .X(_05677_));
 sky130_fd_sc_hd__buf_1 _11456_ (.A(_05677_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_2 _11457_ (.A0(_05639_),
    .A1(net380),
    .S(_05668_),
    .X(_05678_));
 sky130_fd_sc_hd__buf_1 _11458_ (.A(_05678_),
    .X(_00427_));
 sky130_fd_sc_hd__inv_2 _11459_ (.A(net59),
    .Y(_05679_));
 sky130_fd_sc_hd__o21ai_2 _11460_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05643_),
    .Y(_05680_));
 sky130_fd_sc_hd__o21ai_2 _11461_ (.A1(_05679_),
    .A2(_05643_),
    .B1(_05680_),
    .Y(_00428_));
 sky130_fd_sc_hd__and4b_2 _11462_ (.A_N(_04916_),
    .B(_04918_),
    .C(_04920_),
    .D(_04922_),
    .X(_05681_));
 sky130_fd_sc_hd__nor2_2 _11463_ (.A(net136),
    .B(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__a21oi_2 _11464_ (.A1(_05314_),
    .A2(_05681_),
    .B1(_05682_),
    .Y(_00429_));
 sky130_fd_sc_hd__or3_2 _11465_ (.A(_04738_),
    .B(_04739_),
    .C(_05565_),
    .X(_05683_));
 sky130_fd_sc_hd__buf_1 _11466_ (.A(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__mux2_2 _11467_ (.A0(_05318_),
    .A1(net681),
    .S(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__buf_1 _11468_ (.A(_05685_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_2 _11469_ (.A0(_05322_),
    .A1(net253),
    .S(_05684_),
    .X(_05686_));
 sky130_fd_sc_hd__buf_1 _11470_ (.A(_05686_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_2 _11471_ (.A0(_05531_),
    .A1(\rvsingle.dp.rf.rf[12][3] ),
    .S(_05684_),
    .X(_05687_));
 sky130_fd_sc_hd__buf_1 _11472_ (.A(_05687_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_2 _11473_ (.A0(_05377_),
    .A1(net623),
    .S(_05684_),
    .X(_05688_));
 sky130_fd_sc_hd__buf_1 _11474_ (.A(_05688_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_2 _11475_ (.A0(_05534_),
    .A1(\rvsingle.dp.rf.rf[12][5] ),
    .S(_05684_),
    .X(_05689_));
 sky130_fd_sc_hd__buf_1 _11476_ (.A(_05689_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_2 _11477_ (.A0(_05496_),
    .A1(net627),
    .S(_05684_),
    .X(_05690_));
 sky130_fd_sc_hd__buf_1 _11478_ (.A(_05690_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_2 _11479_ (.A0(_05381_),
    .A1(\rvsingle.dp.rf.rf[12][7] ),
    .S(_05684_),
    .X(_05691_));
 sky130_fd_sc_hd__buf_1 _11480_ (.A(_05691_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_2 _11481_ (.A0(_05330_),
    .A1(net686),
    .S(_05684_),
    .X(_05692_));
 sky130_fd_sc_hd__buf_1 _11482_ (.A(_05692_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_2 _11483_ (.A0(_05428_),
    .A1(net467),
    .S(_05684_),
    .X(_05693_));
 sky130_fd_sc_hd__buf_1 _11484_ (.A(_05693_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_2 _11485_ (.A0(_05385_),
    .A1(net653),
    .S(_05684_),
    .X(_05694_));
 sky130_fd_sc_hd__buf_1 _11486_ (.A(_05694_),
    .X(_00439_));
 sky130_fd_sc_hd__buf_1 _11487_ (.A(_05683_),
    .X(_05695_));
 sky130_fd_sc_hd__mux2_2 _11488_ (.A0(_05334_),
    .A1(net566),
    .S(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__buf_1 _11489_ (.A(_05696_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_2 _11490_ (.A0(_04795_),
    .A1(net663),
    .S(_05695_),
    .X(_05697_));
 sky130_fd_sc_hd__buf_1 _11491_ (.A(_05697_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_2 _11492_ (.A0(_04801_),
    .A1(net682),
    .S(_05695_),
    .X(_05698_));
 sky130_fd_sc_hd__buf_1 _11493_ (.A(_05698_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_2 _11494_ (.A0(_05391_),
    .A1(net368),
    .S(_05695_),
    .X(_05699_));
 sky130_fd_sc_hd__buf_1 _11495_ (.A(_05699_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_2 _11496_ (.A0(_04813_),
    .A1(net338),
    .S(_05695_),
    .X(_05700_));
 sky130_fd_sc_hd__buf_1 _11497_ (.A(_05700_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_2 _11498_ (.A0(_05291_),
    .A1(net387),
    .S(_05695_),
    .X(_05701_));
 sky130_fd_sc_hd__buf_1 _11499_ (.A(_05701_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_2 _11500_ (.A0(_05476_),
    .A1(net282),
    .S(_05695_),
    .X(_05702_));
 sky130_fd_sc_hd__buf_1 _11501_ (.A(_05702_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_2 _11502_ (.A0(_05439_),
    .A1(net628),
    .S(_05695_),
    .X(_05703_));
 sky130_fd_sc_hd__buf_1 _11503_ (.A(_05703_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_2 _11504_ (.A0(_05295_),
    .A1(net695),
    .S(_05695_),
    .X(_05704_));
 sky130_fd_sc_hd__buf_1 _11505_ (.A(_05704_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_2 _11506_ (.A0(_05398_),
    .A1(net736),
    .S(_05695_),
    .X(_05705_));
 sky130_fd_sc_hd__buf_1 _11507_ (.A(_05705_),
    .X(_00449_));
 sky130_fd_sc_hd__buf_1 _11508_ (.A(_05683_),
    .X(_05706_));
 sky130_fd_sc_hd__mux2_2 _11509_ (.A0(_05400_),
    .A1(net569),
    .S(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__buf_1 _11510_ (.A(_05707_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_2 _11511_ (.A0(_05300_),
    .A1(\rvsingle.dp.rf.rf[12][22] ),
    .S(_05706_),
    .X(_05708_));
 sky130_fd_sc_hd__buf_1 _11512_ (.A(_05708_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_2 _11513_ (.A0(_05352_),
    .A1(\rvsingle.dp.rf.rf[12][23] ),
    .S(_05706_),
    .X(_05709_));
 sky130_fd_sc_hd__buf_1 _11514_ (.A(_05709_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_2 _11515_ (.A0(_05354_),
    .A1(\rvsingle.dp.rf.rf[12][24] ),
    .S(_05706_),
    .X(_05710_));
 sky130_fd_sc_hd__buf_1 _11516_ (.A(_05710_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_2 _11517_ (.A0(_05304_),
    .A1(net631),
    .S(_05706_),
    .X(_05711_));
 sky130_fd_sc_hd__buf_1 _11518_ (.A(_05711_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_2 _11519_ (.A0(_05407_),
    .A1(net556),
    .S(_05706_),
    .X(_05712_));
 sky130_fd_sc_hd__buf_1 _11520_ (.A(_05712_),
    .X(_00455_));
 sky130_fd_sc_hd__buf_1 _11521_ (.A(_04885_),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_2 _11522_ (.A0(_05713_),
    .A1(net395),
    .S(_05706_),
    .X(_05714_));
 sky130_fd_sc_hd__buf_1 _11523_ (.A(_05714_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_2 _11524_ (.A0(_05359_),
    .A1(net309),
    .S(_05706_),
    .X(_05715_));
 sky130_fd_sc_hd__buf_1 _11525_ (.A(_05715_),
    .X(_00457_));
 sky130_fd_sc_hd__buf_1 _11526_ (.A(_04897_),
    .X(_05716_));
 sky130_fd_sc_hd__mux2_2 _11527_ (.A0(_05716_),
    .A1(net222),
    .S(_05706_),
    .X(_05717_));
 sky130_fd_sc_hd__buf_1 _11528_ (.A(_05717_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_2 _11529_ (.A0(_05639_),
    .A1(net263),
    .S(_05706_),
    .X(_05718_));
 sky130_fd_sc_hd__buf_1 _11530_ (.A(_05718_),
    .X(_00459_));
 sky130_fd_sc_hd__inv_2 _11531_ (.A(net38),
    .Y(_05719_));
 sky130_fd_sc_hd__o21ai_2 _11532_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05681_),
    .Y(_05720_));
 sky130_fd_sc_hd__o21ai_2 _11533_ (.A1(_05719_),
    .A2(_05681_),
    .B1(_05720_),
    .Y(_00460_));
 sky130_fd_sc_hd__buf_1 _11534_ (.A(_04718_),
    .X(_05721_));
 sky130_fd_sc_hd__and4_2 _11535_ (.A(_04720_),
    .B(_05142_),
    .C(_04967_),
    .D(_04968_),
    .X(_05722_));
 sky130_fd_sc_hd__o31a_2 _11536_ (.A1(_04976_),
    .A2(_05417_),
    .A3(_05149_),
    .B1(_02873_),
    .X(_05723_));
 sky130_fd_sc_hd__a21oi_2 _11537_ (.A1(_05721_),
    .A2(_05722_),
    .B1(_05723_),
    .Y(_00461_));
 sky130_fd_sc_hd__buf_1 _11538_ (.A(_04735_),
    .X(_05724_));
 sky130_fd_sc_hd__or3_2 _11539_ (.A(_04976_),
    .B(_04975_),
    .C(_05149_),
    .X(_05725_));
 sky130_fd_sc_hd__buf_1 _11540_ (.A(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__mux2_2 _11541_ (.A0(_05724_),
    .A1(net715),
    .S(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__buf_1 _11542_ (.A(_05727_),
    .X(_00462_));
 sky130_fd_sc_hd__buf_1 _11543_ (.A(_04746_),
    .X(_05728_));
 sky130_fd_sc_hd__buf_1 _11544_ (.A(_05725_),
    .X(_05729_));
 sky130_fd_sc_hd__mux2_2 _11545_ (.A0(_05728_),
    .A1(\rvsingle.dp.rf.rf[11][2] ),
    .S(_05729_),
    .X(_05730_));
 sky130_fd_sc_hd__buf_1 _11546_ (.A(_05730_),
    .X(_00463_));
 sky130_fd_sc_hd__buf_1 _11547_ (.A(_05726_),
    .X(_05731_));
 sky130_fd_sc_hd__buf_1 _11548_ (.A(_04968_),
    .X(_05732_));
 sky130_fd_sc_hd__buf_1 _11549_ (.A(_04967_),
    .X(_05733_));
 sky130_fd_sc_hd__and4_2 _11550_ (.A(_04754_),
    .B(_05732_),
    .C(_05733_),
    .D(_05060_),
    .X(_05734_));
 sky130_fd_sc_hd__a22o_2 _11551_ (.A1(net86),
    .A2(_05731_),
    .B1(_05734_),
    .B2(_05157_),
    .X(_00464_));
 sky130_fd_sc_hd__and4_2 _11552_ (.A(_04759_),
    .B(_05732_),
    .C(_05733_),
    .D(_05060_),
    .X(_05735_));
 sky130_fd_sc_hd__a22o_2 _11553_ (.A1(net113),
    .A2(_05731_),
    .B1(_05735_),
    .B2(_05157_),
    .X(_00465_));
 sky130_fd_sc_hd__and4_2 _11554_ (.A(_04764_),
    .B(_05732_),
    .C(_05733_),
    .D(_05060_),
    .X(_05736_));
 sky130_fd_sc_hd__buf_1 _11555_ (.A(_05146_),
    .X(_05737_));
 sky130_fd_sc_hd__a22o_2 _11556_ (.A1(net125),
    .A2(_05731_),
    .B1(_05736_),
    .B2(_05737_),
    .X(_00466_));
 sky130_fd_sc_hd__and4_2 _11557_ (.A(_04769_),
    .B(_05732_),
    .C(_05733_),
    .D(_05097_),
    .X(_05738_));
 sky130_fd_sc_hd__a22o_2 _11558_ (.A1(net60),
    .A2(_05731_),
    .B1(_05738_),
    .B2(_05737_),
    .X(_00467_));
 sky130_fd_sc_hd__and4_2 _11559_ (.A(_04773_),
    .B(_05732_),
    .C(_05733_),
    .D(_05097_),
    .X(_05739_));
 sky130_fd_sc_hd__a22o_2 _11560_ (.A1(net11),
    .A2(_05726_),
    .B1(_05739_),
    .B2(_05737_),
    .X(_00468_));
 sky130_fd_sc_hd__buf_1 _11561_ (.A(_04777_),
    .X(_05740_));
 sky130_fd_sc_hd__mux2_2 _11562_ (.A0(_05740_),
    .A1(\rvsingle.dp.rf.rf[11][8] ),
    .S(_05729_),
    .X(_05741_));
 sky130_fd_sc_hd__buf_1 _11563_ (.A(_05741_),
    .X(_00469_));
 sky130_fd_sc_hd__and4_2 _11564_ (.A(_04781_),
    .B(_05732_),
    .C(_05733_),
    .D(_05097_),
    .X(_05742_));
 sky130_fd_sc_hd__a22o_2 _11565_ (.A1(net14),
    .A2(_05726_),
    .B1(_05742_),
    .B2(_05737_),
    .X(_00470_));
 sky130_fd_sc_hd__and4_2 _11566_ (.A(_04785_),
    .B(_05732_),
    .C(_05733_),
    .D(_05060_),
    .X(_05743_));
 sky130_fd_sc_hd__a22o_2 _11567_ (.A1(net93),
    .A2(_05726_),
    .B1(_05743_),
    .B2(_05737_),
    .X(_00471_));
 sky130_fd_sc_hd__buf_1 _11568_ (.A(_04789_),
    .X(_05744_));
 sky130_fd_sc_hd__and4_2 _11569_ (.A(_05744_),
    .B(_05732_),
    .C(_05733_),
    .D(_05097_),
    .X(_05745_));
 sky130_fd_sc_hd__a22o_2 _11570_ (.A1(net160),
    .A2(_05726_),
    .B1(_05745_),
    .B2(_05737_),
    .X(_00472_));
 sky130_fd_sc_hd__nand2_2 _11571_ (.A(_04796_),
    .B(_04973_),
    .Y(_05746_));
 sky130_fd_sc_hd__a2bb2o_2 _11572_ (.A1_N(_05167_),
    .A2_N(_05746_),
    .B1(_05731_),
    .B2(net143),
    .X(_00473_));
 sky130_fd_sc_hd__nand2_2 _11573_ (.A(_04802_),
    .B(_04973_),
    .Y(_05747_));
 sky130_fd_sc_hd__a2bb2o_2 _11574_ (.A1_N(_05167_),
    .A2_N(_05747_),
    .B1(_05731_),
    .B2(net157),
    .X(_00474_));
 sky130_fd_sc_hd__or3b_2 _11575_ (.A(_04976_),
    .B(_05417_),
    .C_N(_04807_),
    .X(_05748_));
 sky130_fd_sc_hd__a2bb2o_2 _11576_ (.A1_N(_05167_),
    .A2_N(_05748_),
    .B1(_05731_),
    .B2(net172),
    .X(_00475_));
 sky130_fd_sc_hd__nand2_2 _11577_ (.A(_04814_),
    .B(_04973_),
    .Y(_05749_));
 sky130_fd_sc_hd__a2bb2o_2 _11578_ (.A1_N(_05167_),
    .A2_N(_05749_),
    .B1(_05731_),
    .B2(net104),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_2 _11579_ (.A0(_05344_),
    .A1(net690),
    .S(_05729_),
    .X(_05750_));
 sky130_fd_sc_hd__buf_1 _11580_ (.A(_05750_),
    .X(_00477_));
 sky130_fd_sc_hd__and4_2 _11581_ (.A(_04823_),
    .B(_05732_),
    .C(_05733_),
    .D(_05097_),
    .X(_05751_));
 sky130_fd_sc_hd__a22o_2 _11582_ (.A1(net163),
    .A2(_05726_),
    .B1(_05751_),
    .B2(_05737_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_2 _11583_ (.A0(_05439_),
    .A1(net541),
    .S(_05729_),
    .X(_05752_));
 sky130_fd_sc_hd__buf_1 _11584_ (.A(_05752_),
    .X(_00479_));
 sky130_fd_sc_hd__nand2_2 _11585_ (.A(_04834_),
    .B(_04972_),
    .Y(_05753_));
 sky130_fd_sc_hd__a2bb2o_2 _11586_ (.A1_N(_05167_),
    .A2_N(_05753_),
    .B1(_05731_),
    .B2(net175),
    .X(_00480_));
 sky130_fd_sc_hd__and4_2 _11587_ (.A(_04839_),
    .B(_05732_),
    .C(_05733_),
    .D(_05060_),
    .X(_05754_));
 sky130_fd_sc_hd__a22o_2 _11588_ (.A1(net31),
    .A2(_05726_),
    .B1(_05754_),
    .B2(_05737_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_2 _11589_ (.A0(_05400_),
    .A1(\rvsingle.dp.rf.rf[11][21] ),
    .S(_05729_),
    .X(_05755_));
 sky130_fd_sc_hd__buf_1 _11590_ (.A(_05755_),
    .X(_00482_));
 sky130_fd_sc_hd__and4_2 _11591_ (.A(_04852_),
    .B(_04968_),
    .C(_04967_),
    .D(_05097_),
    .X(_05756_));
 sky130_fd_sc_hd__a22o_2 _11592_ (.A1(net76),
    .A2(_05726_),
    .B1(_05756_),
    .B2(_05737_),
    .X(_00483_));
 sky130_fd_sc_hd__buf_1 _11593_ (.A(_04858_),
    .X(_05757_));
 sky130_fd_sc_hd__mux2_2 _11594_ (.A0(_05757_),
    .A1(net486),
    .S(_05729_),
    .X(_05758_));
 sky130_fd_sc_hd__buf_1 _11595_ (.A(_05758_),
    .X(_00484_));
 sky130_fd_sc_hd__nand2_2 _11596_ (.A(_04863_),
    .B(_04973_),
    .Y(_05759_));
 sky130_fd_sc_hd__a2bb2o_2 _11597_ (.A1_N(_05149_),
    .A2_N(_05759_),
    .B1(_05731_),
    .B2(net102),
    .X(_00485_));
 sky130_fd_sc_hd__and4_2 _11598_ (.A(_04869_),
    .B(_04968_),
    .C(_04967_),
    .D(_05097_),
    .X(_05760_));
 sky130_fd_sc_hd__a22o_2 _11599_ (.A1(net185),
    .A2(_05726_),
    .B1(_05760_),
    .B2(_05737_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_2 _11600_ (.A0(_05407_),
    .A1(net617),
    .S(_05729_),
    .X(_05761_));
 sky130_fd_sc_hd__buf_1 _11601_ (.A(_05761_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_2 _11602_ (.A0(_05713_),
    .A1(net299),
    .S(_05729_),
    .X(_05762_));
 sky130_fd_sc_hd__buf_1 _11603_ (.A(_05762_),
    .X(_00488_));
 sky130_fd_sc_hd__buf_1 _11604_ (.A(_04891_),
    .X(_05763_));
 sky130_fd_sc_hd__mux2_2 _11605_ (.A0(_05763_),
    .A1(net442),
    .S(_05729_),
    .X(_05764_));
 sky130_fd_sc_hd__buf_1 _11606_ (.A(_05764_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_2 _11607_ (.A0(_05716_),
    .A1(net255),
    .S(_05729_),
    .X(_05765_));
 sky130_fd_sc_hd__buf_1 _11608_ (.A(_05765_),
    .X(_00490_));
 sky130_fd_sc_hd__buf_1 _11609_ (.A(_04972_),
    .X(_05766_));
 sky130_fd_sc_hd__o31a_2 _11610_ (.A1(_04976_),
    .A2(_05417_),
    .A3(_05149_),
    .B1(net564),
    .X(_05767_));
 sky130_fd_sc_hd__a31o_2 _11611_ (.A1(_04904_),
    .A2(_05766_),
    .A3(_05146_),
    .B1(_05767_),
    .X(_00491_));
 sky130_fd_sc_hd__inv_2 _11612_ (.A(net55),
    .Y(_05768_));
 sky130_fd_sc_hd__buf_1 _11613_ (.A(_04908_),
    .X(_05769_));
 sky130_fd_sc_hd__buf_1 _11614_ (.A(_04912_),
    .X(_05770_));
 sky130_fd_sc_hd__o21ai_2 _11615_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05722_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21ai_2 _11616_ (.A1(_05768_),
    .A2(_05722_),
    .B1(_05771_),
    .Y(_00492_));
 sky130_fd_sc_hd__and4_2 _11617_ (.A(_04720_),
    .B(_05367_),
    .C(_04967_),
    .D(_04968_),
    .X(_05772_));
 sky130_fd_sc_hd__a21oi_2 _11618_ (.A1(_04973_),
    .A2(_05457_),
    .B1(net109),
    .Y(_05773_));
 sky130_fd_sc_hd__a21oi_2 _11619_ (.A1(_05721_),
    .A2(_05772_),
    .B1(_05773_),
    .Y(_00493_));
 sky130_fd_sc_hd__or3_2 _11620_ (.A(_04976_),
    .B(_05417_),
    .C(_05371_),
    .X(_05774_));
 sky130_fd_sc_hd__buf_1 _11621_ (.A(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__mux2_2 _11622_ (.A0(_05724_),
    .A1(net563),
    .S(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__buf_1 _11623_ (.A(_05776_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_2 _11624_ (.A0(_05728_),
    .A1(net483),
    .S(_05775_),
    .X(_05777_));
 sky130_fd_sc_hd__buf_1 _11625_ (.A(_05777_),
    .X(_00495_));
 sky130_fd_sc_hd__buf_1 _11626_ (.A(_05774_),
    .X(_05778_));
 sky130_fd_sc_hd__buf_1 _11627_ (.A(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__a22o_2 _11628_ (.A1(net204),
    .A2(_05779_),
    .B1(_05734_),
    .B2(_05501_),
    .X(_00496_));
 sky130_fd_sc_hd__a22o_2 _11629_ (.A1(net140),
    .A2(_05779_),
    .B1(_05735_),
    .B2(_05501_),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_2 _11630_ (.A1(net196),
    .A2(_05779_),
    .B1(_05736_),
    .B2(_05501_),
    .X(_00498_));
 sky130_fd_sc_hd__a22o_2 _11631_ (.A1(net63),
    .A2(_05778_),
    .B1(_05738_),
    .B2(_05501_),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_2 _11632_ (.A1(net72),
    .A2(_05778_),
    .B1(_05739_),
    .B2(_05501_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_2 _11633_ (.A0(_05740_),
    .A1(net332),
    .S(_05775_),
    .X(_05780_));
 sky130_fd_sc_hd__buf_1 _11634_ (.A(_05780_),
    .X(_00501_));
 sky130_fd_sc_hd__a22o_2 _11635_ (.A1(net107),
    .A2(_05778_),
    .B1(_05742_),
    .B2(_05501_),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_2 _11636_ (.A1(net18),
    .A2(_05778_),
    .B1(_05743_),
    .B2(_05501_),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_2 _11637_ (.A1(net189),
    .A2(_05778_),
    .B1(_05745_),
    .B2(_05501_),
    .X(_00504_));
 sky130_fd_sc_hd__a2bb2o_2 _11638_ (.A1_N(_05471_),
    .A2_N(_05746_),
    .B1(_05779_),
    .B2(net87),
    .X(_00505_));
 sky130_fd_sc_hd__a2bb2o_2 _11639_ (.A1_N(_05471_),
    .A2_N(_05747_),
    .B1(_05779_),
    .B2(net131),
    .X(_00506_));
 sky130_fd_sc_hd__a2bb2o_2 _11640_ (.A1_N(_05471_),
    .A2_N(_05748_),
    .B1(_05779_),
    .B2(net126),
    .X(_00507_));
 sky130_fd_sc_hd__a2bb2o_2 _11641_ (.A1_N(_05471_),
    .A2_N(_05749_),
    .B1(_05779_),
    .B2(net202),
    .X(_00508_));
 sky130_fd_sc_hd__nand2_2 _11642_ (.A(_04818_),
    .B(_04973_),
    .Y(_05781_));
 sky130_fd_sc_hd__a2bb2o_2 _11643_ (.A1_N(_05471_),
    .A2_N(_05781_),
    .B1(_05779_),
    .B2(net217),
    .X(_00509_));
 sky130_fd_sc_hd__a22o_2 _11644_ (.A1(net199),
    .A2(_05778_),
    .B1(_05751_),
    .B2(_05457_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_2 _11645_ (.A0(_05439_),
    .A1(\rvsingle.dp.rf.rf[19][18] ),
    .S(_05775_),
    .X(_05782_));
 sky130_fd_sc_hd__buf_1 _11646_ (.A(_05782_),
    .X(_00511_));
 sky130_fd_sc_hd__a2bb2o_2 _11647_ (.A1_N(_05371_),
    .A2_N(_05753_),
    .B1(_05779_),
    .B2(net133),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_2 _11648_ (.A1(net65),
    .A2(_05778_),
    .B1(_05754_),
    .B2(_05457_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_2 _11649_ (.A0(_05400_),
    .A1(net813),
    .S(_05775_),
    .X(_05783_));
 sky130_fd_sc_hd__buf_1 _11650_ (.A(_05783_),
    .X(_00514_));
 sky130_fd_sc_hd__a22o_2 _11651_ (.A1(net200),
    .A2(_05778_),
    .B1(_05756_),
    .B2(_05457_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_2 _11652_ (.A0(_05757_),
    .A1(net250),
    .S(_05775_),
    .X(_05784_));
 sky130_fd_sc_hd__buf_1 _11653_ (.A(_05784_),
    .X(_00516_));
 sky130_fd_sc_hd__a2bb2o_2 _11654_ (.A1_N(_05371_),
    .A2_N(_05759_),
    .B1(_05779_),
    .B2(net173),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_2 _11655_ (.A1(net213),
    .A2(_05778_),
    .B1(_05760_),
    .B2(_05457_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_2 _11656_ (.A0(_05407_),
    .A1(\rvsingle.dp.rf.rf[19][26] ),
    .S(_05775_),
    .X(_05785_));
 sky130_fd_sc_hd__buf_1 _11657_ (.A(_05785_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_2 _11658_ (.A0(_05713_),
    .A1(net441),
    .S(_05775_),
    .X(_05786_));
 sky130_fd_sc_hd__buf_1 _11659_ (.A(_05786_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_2 _11660_ (.A0(_05763_),
    .A1(net257),
    .S(_05775_),
    .X(_05787_));
 sky130_fd_sc_hd__buf_1 _11661_ (.A(_05787_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_2 _11662_ (.A0(_05716_),
    .A1(net285),
    .S(_05775_),
    .X(_05788_));
 sky130_fd_sc_hd__buf_1 _11663_ (.A(_05788_),
    .X(_00522_));
 sky130_fd_sc_hd__o31a_2 _11664_ (.A1(_04976_),
    .A2(_05417_),
    .A3(_05371_),
    .B1(net518),
    .X(_05789_));
 sky130_fd_sc_hd__a31o_2 _11665_ (.A1(_04904_),
    .A2(_05766_),
    .A3(_05457_),
    .B1(_05789_),
    .X(_00523_));
 sky130_fd_sc_hd__inv_2 _11666_ (.A(net51),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ai_2 _11667_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05772_),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_2 _11668_ (.A1(_05790_),
    .A2(_05772_),
    .B1(_05791_),
    .Y(_00524_));
 sky130_fd_sc_hd__and3_2 _11669_ (.A(_04720_),
    .B(_04728_),
    .C(_05142_),
    .X(_05792_));
 sky130_fd_sc_hd__nor2_2 _11670_ (.A(net187),
    .B(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__a21oi_2 _11671_ (.A1(_05721_),
    .A2(_05792_),
    .B1(_05793_),
    .Y(_00525_));
 sky130_fd_sc_hd__or4b_2 _11672_ (.A(_04738_),
    .B(_04733_),
    .C(_05149_),
    .D_N(_04739_),
    .X(_05794_));
 sky130_fd_sc_hd__buf_1 _11673_ (.A(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__mux2_2 _11674_ (.A0(_05724_),
    .A1(\rvsingle.dp.rf.rf[10][1] ),
    .S(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__buf_1 _11675_ (.A(_05796_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_2 _11676_ (.A0(_05728_),
    .A1(\rvsingle.dp.rf.rf[10][2] ),
    .S(_05795_),
    .X(_05797_));
 sky130_fd_sc_hd__buf_1 _11677_ (.A(_05797_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_2 _11678_ (.A0(_05531_),
    .A1(\rvsingle.dp.rf.rf[10][3] ),
    .S(_05795_),
    .X(_05798_));
 sky130_fd_sc_hd__buf_1 _11679_ (.A(_05798_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_2 _11680_ (.A0(_05377_),
    .A1(net598),
    .S(_05795_),
    .X(_05799_));
 sky130_fd_sc_hd__buf_1 _11681_ (.A(_05799_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_2 _11682_ (.A0(_05534_),
    .A1(\rvsingle.dp.rf.rf[10][5] ),
    .S(_05795_),
    .X(_05800_));
 sky130_fd_sc_hd__buf_1 _11683_ (.A(_05800_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_2 _11684_ (.A0(_05496_),
    .A1(net719),
    .S(_05795_),
    .X(_05801_));
 sky130_fd_sc_hd__buf_1 _11685_ (.A(_05801_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_2 _11686_ (.A0(_05381_),
    .A1(\rvsingle.dp.rf.rf[10][7] ),
    .S(_05795_),
    .X(_05802_));
 sky130_fd_sc_hd__buf_1 _11687_ (.A(_05802_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_2 _11688_ (.A0(_05740_),
    .A1(net632),
    .S(_05795_),
    .X(_05803_));
 sky130_fd_sc_hd__buf_1 _11689_ (.A(_05803_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_2 _11690_ (.A0(_05428_),
    .A1(net397),
    .S(_05795_),
    .X(_05804_));
 sky130_fd_sc_hd__buf_1 _11691_ (.A(_05804_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_2 _11692_ (.A0(_05385_),
    .A1(net516),
    .S(_05795_),
    .X(_05805_));
 sky130_fd_sc_hd__buf_1 _11693_ (.A(_05805_),
    .X(_00535_));
 sky130_fd_sc_hd__buf_1 _11694_ (.A(_05794_),
    .X(_05806_));
 sky130_fd_sc_hd__mux2_2 _11695_ (.A0(_05744_),
    .A1(\rvsingle.dp.rf.rf[10][11] ),
    .S(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__buf_1 _11696_ (.A(_05807_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_2 _11697_ (.A0(_04795_),
    .A1(net363),
    .S(_05806_),
    .X(_05808_));
 sky130_fd_sc_hd__buf_1 _11698_ (.A(_05808_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_2 _11699_ (.A0(_04801_),
    .A1(net493),
    .S(_05806_),
    .X(_05809_));
 sky130_fd_sc_hd__buf_1 _11700_ (.A(_05809_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_2 _11701_ (.A0(_05391_),
    .A1(\rvsingle.dp.rf.rf[10][14] ),
    .S(_05806_),
    .X(_05810_));
 sky130_fd_sc_hd__buf_1 _11702_ (.A(_05810_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_2 _11703_ (.A0(_04813_),
    .A1(net552),
    .S(_05806_),
    .X(_05811_));
 sky130_fd_sc_hd__buf_1 _11704_ (.A(_05811_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_2 _11705_ (.A0(_05344_),
    .A1(net346),
    .S(_05806_),
    .X(_05812_));
 sky130_fd_sc_hd__buf_1 _11706_ (.A(_05812_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_2 _11707_ (.A0(_05476_),
    .A1(\rvsingle.dp.rf.rf[10][17] ),
    .S(_05806_),
    .X(_05813_));
 sky130_fd_sc_hd__buf_1 _11708_ (.A(_05813_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_2 _11709_ (.A0(_05439_),
    .A1(net412),
    .S(_05806_),
    .X(_05814_));
 sky130_fd_sc_hd__buf_1 _11710_ (.A(_05814_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_2 _11711_ (.A0(_05295_),
    .A1(\rvsingle.dp.rf.rf[10][19] ),
    .S(_05806_),
    .X(_05815_));
 sky130_fd_sc_hd__buf_1 _11712_ (.A(_05815_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_2 _11713_ (.A0(_05398_),
    .A1(\rvsingle.dp.rf.rf[10][20] ),
    .S(_05806_),
    .X(_05816_));
 sky130_fd_sc_hd__buf_1 _11714_ (.A(_05816_),
    .X(_00545_));
 sky130_fd_sc_hd__buf_1 _11715_ (.A(_05794_),
    .X(_05817_));
 sky130_fd_sc_hd__mux2_2 _11716_ (.A0(_04845_),
    .A1(net422),
    .S(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__buf_1 _11717_ (.A(_05818_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_2 _11718_ (.A0(_05300_),
    .A1(net587),
    .S(_05817_),
    .X(_05819_));
 sky130_fd_sc_hd__buf_1 _11719_ (.A(_05819_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_2 _11720_ (.A0(_05757_),
    .A1(net584),
    .S(_05817_),
    .X(_05820_));
 sky130_fd_sc_hd__buf_1 _11721_ (.A(_05820_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_2 _11722_ (.A0(_05354_),
    .A1(net259),
    .S(_05817_),
    .X(_05821_));
 sky130_fd_sc_hd__buf_1 _11723_ (.A(_05821_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_2 _11724_ (.A0(_05304_),
    .A1(net743),
    .S(_05817_),
    .X(_05822_));
 sky130_fd_sc_hd__buf_1 _11725_ (.A(_05822_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_2 _11726_ (.A0(_04876_),
    .A1(net550),
    .S(_05817_),
    .X(_05823_));
 sky130_fd_sc_hd__buf_1 _11727_ (.A(_05823_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_2 _11728_ (.A0(_05713_),
    .A1(net379),
    .S(_05817_),
    .X(_05824_));
 sky130_fd_sc_hd__buf_1 _11729_ (.A(_05824_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_2 _11730_ (.A0(_05763_),
    .A1(net281),
    .S(_05817_),
    .X(_05825_));
 sky130_fd_sc_hd__buf_1 _11731_ (.A(_05825_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_2 _11732_ (.A0(_05716_),
    .A1(net287),
    .S(_05817_),
    .X(_05826_));
 sky130_fd_sc_hd__buf_1 _11733_ (.A(_05826_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_2 _11734_ (.A0(_05639_),
    .A1(net452),
    .S(_05817_),
    .X(_05827_));
 sky130_fd_sc_hd__buf_1 _11735_ (.A(_05827_),
    .X(_00555_));
 sky130_fd_sc_hd__inv_2 _11736_ (.A(net48),
    .Y(_05828_));
 sky130_fd_sc_hd__o21ai_2 _11737_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05792_),
    .Y(_05829_));
 sky130_fd_sc_hd__o21ai_2 _11738_ (.A1(_05828_),
    .A2(_05792_),
    .B1(_05829_),
    .Y(_00556_));
 sky130_fd_sc_hd__nor3b_2 _11739_ (.A(_04915_),
    .B(_04917_),
    .C_N(_04965_),
    .Y(_05830_));
 sky130_fd_sc_hd__and4_2 _11740_ (.A(_04720_),
    .B(_05830_),
    .C(_04967_),
    .D(_04968_),
    .X(_05831_));
 sky130_fd_sc_hd__buf_1 _11741_ (.A(_05830_),
    .X(_05832_));
 sky130_fd_sc_hd__a21oi_2 _11742_ (.A1(_04973_),
    .A2(_05832_),
    .B1(net79),
    .Y(_05833_));
 sky130_fd_sc_hd__a21oi_2 _11743_ (.A1(_05721_),
    .A2(_05831_),
    .B1(_05833_),
    .Y(_00557_));
 sky130_fd_sc_hd__or3b_2 _11744_ (.A(_04722_),
    .B(_04723_),
    .C_N(_04724_),
    .X(_05834_));
 sky130_fd_sc_hd__buf_1 _11745_ (.A(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__a311o_2 _11746_ (.A1(_04505_),
    .A2(_01071_),
    .A3(_01062_),
    .B1(_05417_),
    .C1(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__buf_1 _11747_ (.A(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__mux2_2 _11748_ (.A0(_05724_),
    .A1(net808),
    .S(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__buf_1 _11749_ (.A(_05838_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_2 _11750_ (.A0(_05728_),
    .A1(net799),
    .S(_05837_),
    .X(_05839_));
 sky130_fd_sc_hd__buf_1 _11751_ (.A(_05839_),
    .X(_00559_));
 sky130_fd_sc_hd__buf_1 _11752_ (.A(_05837_),
    .X(_05840_));
 sky130_fd_sc_hd__buf_1 _11753_ (.A(_05830_),
    .X(_05841_));
 sky130_fd_sc_hd__a22o_2 _11754_ (.A1(_05840_),
    .A2(net37),
    .B1(_05734_),
    .B2(_05841_),
    .X(_00560_));
 sky130_fd_sc_hd__a22o_2 _11755_ (.A1(_05840_),
    .A2(net36),
    .B1(_05735_),
    .B2(_05841_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_2 _11756_ (.A0(_05534_),
    .A1(\rvsingle.dp.rf.rf[7][5] ),
    .S(_05837_),
    .X(_05842_));
 sky130_fd_sc_hd__buf_1 _11757_ (.A(_05842_),
    .X(_00562_));
 sky130_fd_sc_hd__a22o_2 _11758_ (.A1(_05840_),
    .A2(net117),
    .B1(_05738_),
    .B2(_05841_),
    .X(_00563_));
 sky130_fd_sc_hd__a22o_2 _11759_ (.A1(_05840_),
    .A2(net92),
    .B1(_05739_),
    .B2(_05841_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_2 _11760_ (.A0(_05740_),
    .A1(net649),
    .S(_05837_),
    .X(_05843_));
 sky130_fd_sc_hd__buf_1 _11761_ (.A(_05843_),
    .X(_00565_));
 sky130_fd_sc_hd__a22o_2 _11762_ (.A1(_05840_),
    .A2(net91),
    .B1(_05742_),
    .B2(_05841_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_2 _11763_ (.A0(_05385_),
    .A1(net588),
    .S(_05837_),
    .X(_05844_));
 sky130_fd_sc_hd__buf_1 _11764_ (.A(_05844_),
    .X(_00567_));
 sky130_fd_sc_hd__a22o_2 _11765_ (.A1(_05837_),
    .A2(net101),
    .B1(_05745_),
    .B2(_05841_),
    .X(_00568_));
 sky130_fd_sc_hd__buf_1 _11766_ (.A(_05836_),
    .X(_05845_));
 sky130_fd_sc_hd__mux2_2 _11767_ (.A0(_04795_),
    .A1(net251),
    .S(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__buf_1 _11768_ (.A(_05846_),
    .X(_00569_));
 sky130_fd_sc_hd__buf_1 _11769_ (.A(_05835_),
    .X(_05847_));
 sky130_fd_sc_hd__a2bb2o_2 _11770_ (.A1_N(_05747_),
    .A2_N(_05847_),
    .B1(_05840_),
    .B2(net165),
    .X(_00570_));
 sky130_fd_sc_hd__a2bb2o_2 _11771_ (.A1_N(_05748_),
    .A2_N(_05847_),
    .B1(_05840_),
    .B2(net95),
    .X(_00571_));
 sky130_fd_sc_hd__a2bb2o_2 _11772_ (.A1_N(_05749_),
    .A2_N(_05847_),
    .B1(_05840_),
    .B2(net69),
    .X(_00572_));
 sky130_fd_sc_hd__a2bb2o_2 _11773_ (.A1_N(_05781_),
    .A2_N(_05847_),
    .B1(_05840_),
    .B2(net153),
    .X(_00573_));
 sky130_fd_sc_hd__a22o_2 _11774_ (.A1(_05837_),
    .A2(net209),
    .B1(_05751_),
    .B2(_05841_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_2 _11775_ (.A0(_05173_),
    .A1(net714),
    .S(_05845_),
    .X(_05848_));
 sky130_fd_sc_hd__buf_1 _11776_ (.A(_05848_),
    .X(_00575_));
 sky130_fd_sc_hd__a2bb2o_2 _11777_ (.A1_N(_05753_),
    .A2_N(_05847_),
    .B1(_05840_),
    .B2(net105),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_2 _11778_ (.A0(_05398_),
    .A1(net547),
    .S(_05845_),
    .X(_05849_));
 sky130_fd_sc_hd__buf_1 _11779_ (.A(_05849_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_2 _11780_ (.A0(_04845_),
    .A1(net310),
    .S(_05845_),
    .X(_05850_));
 sky130_fd_sc_hd__buf_1 _11781_ (.A(_05850_),
    .X(_00578_));
 sky130_fd_sc_hd__a22o_2 _11782_ (.A1(_05837_),
    .A2(net119),
    .B1(_05756_),
    .B2(_05841_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_2 _11783_ (.A0(_05757_),
    .A1(\rvsingle.dp.rf.rf[7][23] ),
    .S(_05845_),
    .X(_05851_));
 sky130_fd_sc_hd__buf_1 _11784_ (.A(_05851_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_2 _11785_ (.A0(_05132_),
    .A1(net352),
    .S(_05845_),
    .X(_05852_));
 sky130_fd_sc_hd__buf_1 _11786_ (.A(_05852_),
    .X(_00581_));
 sky130_fd_sc_hd__a22o_2 _11787_ (.A1(_05837_),
    .A2(net190),
    .B1(_05760_),
    .B2(_05841_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_2 _11788_ (.A0(_04876_),
    .A1(net660),
    .S(_05845_),
    .X(_05853_));
 sky130_fd_sc_hd__buf_1 _11789_ (.A(_05853_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_2 _11790_ (.A0(_05713_),
    .A1(net497),
    .S(_05845_),
    .X(_05854_));
 sky130_fd_sc_hd__buf_1 _11791_ (.A(_05854_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_2 _11792_ (.A0(_05763_),
    .A1(net277),
    .S(_05845_),
    .X(_05855_));
 sky130_fd_sc_hd__buf_1 _11793_ (.A(_05855_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_2 _11794_ (.A0(_05716_),
    .A1(net359),
    .S(_05845_),
    .X(_05856_));
 sky130_fd_sc_hd__buf_1 _11795_ (.A(_05856_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_2 _11796_ (.A0(_05639_),
    .A1(net699),
    .S(_05836_),
    .X(_05857_));
 sky130_fd_sc_hd__buf_1 _11797_ (.A(_05857_),
    .X(_00587_));
 sky130_fd_sc_hd__inv_2 _11798_ (.A(net32),
    .Y(_05858_));
 sky130_fd_sc_hd__o21ai_2 _11799_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05831_),
    .Y(_05859_));
 sky130_fd_sc_hd__o21ai_2 _11800_ (.A1(_05858_),
    .A2(_05831_),
    .B1(_05859_),
    .Y(_00588_));
 sky130_fd_sc_hd__nor4b_2 _11801_ (.A(_04918_),
    .B(_04928_),
    .C(_05417_),
    .D_N(_04915_),
    .Y(_05860_));
 sky130_fd_sc_hd__nor2_2 _11802_ (.A(net120),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__a21oi_2 _11803_ (.A1(_05721_),
    .A2(_05860_),
    .B1(_05861_),
    .Y(_00589_));
 sky130_fd_sc_hd__or4b_2 _11804_ (.A(_04723_),
    .B(_04928_),
    .C(_04975_),
    .D_N(_04722_),
    .X(_05862_));
 sky130_fd_sc_hd__buf_1 _11805_ (.A(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__mux2_2 _11806_ (.A0(_05724_),
    .A1(net298),
    .S(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__buf_1 _11807_ (.A(_05864_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_2 _11808_ (.A0(_05728_),
    .A1(net721),
    .S(_05863_),
    .X(_05865_));
 sky130_fd_sc_hd__buf_1 _11809_ (.A(_05865_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_2 _11810_ (.A0(_05531_),
    .A1(net758),
    .S(_05863_),
    .X(_05866_));
 sky130_fd_sc_hd__buf_1 _11811_ (.A(_05866_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_2 _11812_ (.A0(_05377_),
    .A1(\rvsingle.dp.rf.rf[23][4] ),
    .S(_05863_),
    .X(_05867_));
 sky130_fd_sc_hd__buf_1 _11813_ (.A(_05867_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_2 _11814_ (.A0(_05534_),
    .A1(net392),
    .S(_05863_),
    .X(_05868_));
 sky130_fd_sc_hd__buf_1 _11815_ (.A(_05868_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_2 _11816_ (.A0(_05496_),
    .A1(net779),
    .S(_05863_),
    .X(_05869_));
 sky130_fd_sc_hd__buf_1 _11817_ (.A(_05869_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_2 _11818_ (.A0(_05381_),
    .A1(net778),
    .S(_05863_),
    .X(_05870_));
 sky130_fd_sc_hd__buf_1 _11819_ (.A(_05870_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_2 _11820_ (.A0(_05740_),
    .A1(net270),
    .S(_05863_),
    .X(_05871_));
 sky130_fd_sc_hd__buf_1 _11821_ (.A(_05871_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_2 _11822_ (.A0(_05428_),
    .A1(net269),
    .S(_05863_),
    .X(_05872_));
 sky130_fd_sc_hd__buf_1 _11823_ (.A(_05872_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_2 _11824_ (.A0(_04785_),
    .A1(net317),
    .S(_05863_),
    .X(_05873_));
 sky130_fd_sc_hd__buf_1 _11825_ (.A(_05873_),
    .X(_00599_));
 sky130_fd_sc_hd__buf_1 _11826_ (.A(_05862_),
    .X(_05874_));
 sky130_fd_sc_hd__mux2_2 _11827_ (.A0(_05744_),
    .A1(net780),
    .S(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__buf_1 _11828_ (.A(_05875_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_2 _11829_ (.A0(_04795_),
    .A1(net696),
    .S(_05874_),
    .X(_05876_));
 sky130_fd_sc_hd__buf_1 _11830_ (.A(_05876_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_2 _11831_ (.A0(_04801_),
    .A1(net498),
    .S(_05874_),
    .X(_05877_));
 sky130_fd_sc_hd__buf_1 _11832_ (.A(_05877_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_2 _11833_ (.A0(_05391_),
    .A1(net246),
    .S(_05874_),
    .X(_05878_));
 sky130_fd_sc_hd__buf_1 _11834_ (.A(_05878_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_2 _11835_ (.A0(_04813_),
    .A1(net675),
    .S(_05874_),
    .X(_05879_));
 sky130_fd_sc_hd__buf_1 _11836_ (.A(_05879_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_2 _11837_ (.A0(_05344_),
    .A1(net333),
    .S(_05874_),
    .X(_05880_));
 sky130_fd_sc_hd__buf_1 _11838_ (.A(_05880_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_2 _11839_ (.A0(_05476_),
    .A1(net562),
    .S(_05874_),
    .X(_05881_));
 sky130_fd_sc_hd__buf_1 _11840_ (.A(_05881_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_2 _11841_ (.A0(_05173_),
    .A1(\rvsingle.dp.rf.rf[23][18] ),
    .S(_05874_),
    .X(_05882_));
 sky130_fd_sc_hd__buf_1 _11842_ (.A(_05882_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_2 _11843_ (.A0(_04833_),
    .A1(net536),
    .S(_05874_),
    .X(_05883_));
 sky130_fd_sc_hd__buf_1 _11844_ (.A(_05883_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_2 _11845_ (.A0(_04839_),
    .A1(net505),
    .S(_05874_),
    .X(_05884_));
 sky130_fd_sc_hd__buf_1 _11846_ (.A(_05884_),
    .X(_00609_));
 sky130_fd_sc_hd__buf_1 _11847_ (.A(_05862_),
    .X(_05885_));
 sky130_fd_sc_hd__mux2_2 _11848_ (.A0(_04845_),
    .A1(net811),
    .S(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__buf_1 _11849_ (.A(_05886_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_2 _11850_ (.A0(_04852_),
    .A1(net635),
    .S(_05885_),
    .X(_05887_));
 sky130_fd_sc_hd__buf_1 _11851_ (.A(_05887_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_2 _11852_ (.A0(_05757_),
    .A1(net256),
    .S(_05885_),
    .X(_05888_));
 sky130_fd_sc_hd__buf_1 _11853_ (.A(_05888_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_2 _11854_ (.A0(_05132_),
    .A1(net568),
    .S(_05885_),
    .X(_05889_));
 sky130_fd_sc_hd__buf_1 _11855_ (.A(_05889_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_2 _11856_ (.A0(_04869_),
    .A1(net477),
    .S(_05885_),
    .X(_05890_));
 sky130_fd_sc_hd__buf_1 _11857_ (.A(_05890_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_2 _11858_ (.A0(_04876_),
    .A1(net691),
    .S(_05885_),
    .X(_05891_));
 sky130_fd_sc_hd__buf_1 _11859_ (.A(_05891_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_2 _11860_ (.A0(_05713_),
    .A1(net784),
    .S(_05885_),
    .X(_05892_));
 sky130_fd_sc_hd__buf_1 _11861_ (.A(_05892_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_2 _11862_ (.A0(_05763_),
    .A1(net235),
    .S(_05885_),
    .X(_05893_));
 sky130_fd_sc_hd__buf_1 _11863_ (.A(_05893_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_2 _11864_ (.A0(_05716_),
    .A1(net661),
    .S(_05885_),
    .X(_05894_));
 sky130_fd_sc_hd__buf_1 _11865_ (.A(_05894_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_2 _11866_ (.A0(_05639_),
    .A1(net266),
    .S(_05885_),
    .X(_05895_));
 sky130_fd_sc_hd__buf_1 _11867_ (.A(_05895_),
    .X(_00619_));
 sky130_fd_sc_hd__inv_2 _11868_ (.A(net44),
    .Y(_05896_));
 sky130_fd_sc_hd__o21ai_2 _11869_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05860_),
    .Y(_05897_));
 sky130_fd_sc_hd__o21ai_2 _11870_ (.A1(_05896_),
    .A2(_05860_),
    .B1(_05897_),
    .Y(_00620_));
 sky130_fd_sc_hd__buf_1 _11871_ (.A(reset),
    .X(_05898_));
 sky130_fd_sc_hd__inv_2 _11872_ (.A(_05898_),
    .Y(_00000_));
 sky130_fd_sc_hd__inv_2 _11873_ (.A(_05898_),
    .Y(_00001_));
 sky130_fd_sc_hd__and3_2 _11874_ (.A(_04720_),
    .B(_04728_),
    .C(_05830_),
    .X(_05899_));
 sky130_fd_sc_hd__nor2_2 _11875_ (.A(net111),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__a21oi_2 _11876_ (.A1(_05721_),
    .A2(_05899_),
    .B1(_05900_),
    .Y(_00623_));
 sky130_fd_sc_hd__or4b_2 _11877_ (.A(_04738_),
    .B(_04733_),
    .C(_05835_),
    .D_N(_04739_),
    .X(_05901_));
 sky130_fd_sc_hd__buf_1 _11878_ (.A(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__mux2_2 _11879_ (.A0(_05724_),
    .A1(\rvsingle.dp.rf.rf[6][1] ),
    .S(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__buf_1 _11880_ (.A(_05903_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_2 _11881_ (.A0(_05728_),
    .A1(\rvsingle.dp.rf.rf[6][2] ),
    .S(_05902_),
    .X(_05904_));
 sky130_fd_sc_hd__buf_1 _11882_ (.A(_05904_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_2 _11883_ (.A0(_05531_),
    .A1(\rvsingle.dp.rf.rf[6][3] ),
    .S(_05902_),
    .X(_05905_));
 sky130_fd_sc_hd__buf_1 _11884_ (.A(_05905_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_2 _11885_ (.A0(_04759_),
    .A1(net542),
    .S(_05902_),
    .X(_05906_));
 sky130_fd_sc_hd__buf_1 _11886_ (.A(_05906_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_2 _11887_ (.A0(_05534_),
    .A1(net734),
    .S(_05902_),
    .X(_05907_));
 sky130_fd_sc_hd__buf_1 _11888_ (.A(_05907_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_2 _11889_ (.A0(_05496_),
    .A1(\rvsingle.dp.rf.rf[6][6] ),
    .S(_05902_),
    .X(_05908_));
 sky130_fd_sc_hd__buf_1 _11890_ (.A(_05908_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_2 _11891_ (.A0(_04773_),
    .A1(net487),
    .S(_05902_),
    .X(_05909_));
 sky130_fd_sc_hd__buf_1 _11892_ (.A(_05909_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_2 _11893_ (.A0(_05740_),
    .A1(net433),
    .S(_05902_),
    .X(_05910_));
 sky130_fd_sc_hd__buf_1 _11894_ (.A(_05910_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_2 _11895_ (.A0(_05428_),
    .A1(net643),
    .S(_05902_),
    .X(_05911_));
 sky130_fd_sc_hd__buf_1 _11896_ (.A(_05911_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_2 _11897_ (.A0(_04785_),
    .A1(net329),
    .S(_05902_),
    .X(_05912_));
 sky130_fd_sc_hd__buf_1 _11898_ (.A(_05912_),
    .X(_00633_));
 sky130_fd_sc_hd__buf_1 _11899_ (.A(_05901_),
    .X(_05913_));
 sky130_fd_sc_hd__mux2_2 _11900_ (.A0(_05744_),
    .A1(net336),
    .S(_05913_),
    .X(_05914_));
 sky130_fd_sc_hd__buf_1 _11901_ (.A(_05914_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_2 _11902_ (.A0(_04795_),
    .A1(net526),
    .S(_05913_),
    .X(_05915_));
 sky130_fd_sc_hd__buf_1 _11903_ (.A(_05915_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_2 _11904_ (.A0(_04801_),
    .A1(net703),
    .S(_05913_),
    .X(_05916_));
 sky130_fd_sc_hd__buf_1 _11905_ (.A(_05916_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_2 _11906_ (.A0(_04807_),
    .A1(net492),
    .S(_05913_),
    .X(_05917_));
 sky130_fd_sc_hd__buf_1 _11907_ (.A(_05917_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_2 _11908_ (.A0(_04813_),
    .A1(net561),
    .S(_05913_),
    .X(_05918_));
 sky130_fd_sc_hd__buf_1 _11909_ (.A(_05918_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_2 _11910_ (.A0(_05344_),
    .A1(net360),
    .S(_05913_),
    .X(_05919_));
 sky130_fd_sc_hd__buf_1 _11911_ (.A(_05919_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_2 _11912_ (.A0(_05476_),
    .A1(net543),
    .S(_05913_),
    .X(_05920_));
 sky130_fd_sc_hd__buf_1 _11913_ (.A(_05920_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_2 _11914_ (.A0(_05173_),
    .A1(net414),
    .S(_05913_),
    .X(_05921_));
 sky130_fd_sc_hd__buf_1 _11915_ (.A(_05921_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_2 _11916_ (.A0(_04833_),
    .A1(net520),
    .S(_05913_),
    .X(_05922_));
 sky130_fd_sc_hd__buf_1 _11917_ (.A(_05922_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_2 _11918_ (.A0(_04839_),
    .A1(net665),
    .S(_05913_),
    .X(_05923_));
 sky130_fd_sc_hd__buf_1 _11919_ (.A(_05923_),
    .X(_00643_));
 sky130_fd_sc_hd__buf_1 _11920_ (.A(_05901_),
    .X(_05924_));
 sky130_fd_sc_hd__mux2_2 _11921_ (.A0(_04845_),
    .A1(net384),
    .S(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__buf_1 _11922_ (.A(_05925_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_2 _11923_ (.A0(_04852_),
    .A1(net230),
    .S(_05924_),
    .X(_05926_));
 sky130_fd_sc_hd__buf_1 _11924_ (.A(_05926_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_2 _11925_ (.A0(_05757_),
    .A1(\rvsingle.dp.rf.rf[6][23] ),
    .S(_05924_),
    .X(_05927_));
 sky130_fd_sc_hd__buf_1 _11926_ (.A(_05927_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_2 _11927_ (.A0(_05132_),
    .A1(net249),
    .S(_05924_),
    .X(_05928_));
 sky130_fd_sc_hd__buf_1 _11928_ (.A(_05928_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_2 _11929_ (.A0(_04869_),
    .A1(net260),
    .S(_05924_),
    .X(_05929_));
 sky130_fd_sc_hd__buf_1 _11930_ (.A(_05929_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_2 _11931_ (.A0(_04876_),
    .A1(net579),
    .S(_05924_),
    .X(_05930_));
 sky130_fd_sc_hd__buf_1 _11932_ (.A(_05930_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_2 _11933_ (.A0(_05713_),
    .A1(net240),
    .S(_05924_),
    .X(_05931_));
 sky130_fd_sc_hd__buf_1 _11934_ (.A(_05931_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_2 _11935_ (.A0(_05763_),
    .A1(net292),
    .S(_05924_),
    .X(_05932_));
 sky130_fd_sc_hd__buf_1 _11936_ (.A(_05932_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_2 _11937_ (.A0(_05716_),
    .A1(net377),
    .S(_05924_),
    .X(_05933_));
 sky130_fd_sc_hd__buf_1 _11938_ (.A(_05933_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_2 _11939_ (.A0(_05639_),
    .A1(net553),
    .S(_05924_),
    .X(_05934_));
 sky130_fd_sc_hd__buf_1 _11940_ (.A(_05934_),
    .X(_00653_));
 sky130_fd_sc_hd__inv_2 _11941_ (.A(net43),
    .Y(_05935_));
 sky130_fd_sc_hd__o21ai_2 _11942_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05899_),
    .Y(_05936_));
 sky130_fd_sc_hd__o21ai_2 _11943_ (.A1(_05935_),
    .A2(_05899_),
    .B1(_05936_),
    .Y(_00654_));
 sky130_fd_sc_hd__and3_2 _11944_ (.A(_04721_),
    .B(_04920_),
    .C(_05830_),
    .X(_05937_));
 sky130_fd_sc_hd__a21oi_2 _11945_ (.A1(_05099_),
    .A2(_05832_),
    .B1(net116),
    .Y(_05938_));
 sky130_fd_sc_hd__a21oi_2 _11946_ (.A1(_05721_),
    .A2(_05937_),
    .B1(_05938_),
    .Y(_00655_));
 sky130_fd_sc_hd__or4_2 _11947_ (.A(_04737_),
    .B(_04739_),
    .C(_04976_),
    .D(_05835_),
    .X(_05939_));
 sky130_fd_sc_hd__buf_1 _11948_ (.A(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__mux2_2 _11949_ (.A0(_05724_),
    .A1(\rvsingle.dp.rf.rf[4][1] ),
    .S(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__buf_1 _11950_ (.A(_05941_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_2 _11951_ (.A0(_05728_),
    .A1(\rvsingle.dp.rf.rf[4][2] ),
    .S(_05940_),
    .X(_05942_));
 sky130_fd_sc_hd__buf_1 _11952_ (.A(_05942_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_2 _11953_ (.A0(_05531_),
    .A1(\rvsingle.dp.rf.rf[4][3] ),
    .S(_05940_),
    .X(_05943_));
 sky130_fd_sc_hd__buf_1 _11954_ (.A(_05943_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_2 _11955_ (.A0(_04759_),
    .A1(net275),
    .S(_05940_),
    .X(_05944_));
 sky130_fd_sc_hd__buf_1 _11956_ (.A(_05944_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_2 _11957_ (.A0(_05534_),
    .A1(net679),
    .S(_05940_),
    .X(_05945_));
 sky130_fd_sc_hd__buf_1 _11958_ (.A(_05945_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_2 _11959_ (.A0(_05496_),
    .A1(\rvsingle.dp.rf.rf[4][6] ),
    .S(_05940_),
    .X(_05946_));
 sky130_fd_sc_hd__buf_1 _11960_ (.A(_05946_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_2 _11961_ (.A0(_04773_),
    .A1(net549),
    .S(_05940_),
    .X(_05947_));
 sky130_fd_sc_hd__buf_1 _11962_ (.A(_05947_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_2 _11963_ (.A0(_05740_),
    .A1(net314),
    .S(_05940_),
    .X(_05948_));
 sky130_fd_sc_hd__buf_1 _11964_ (.A(_05948_),
    .X(_00663_));
 sky130_fd_sc_hd__buf_1 _11965_ (.A(_05939_),
    .X(_05949_));
 sky130_fd_sc_hd__mux2_2 _11966_ (.A0(_04781_),
    .A1(net751),
    .S(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__buf_1 _11967_ (.A(_05950_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_2 _11968_ (.A0(_04785_),
    .A1(net560),
    .S(_05949_),
    .X(_05951_));
 sky130_fd_sc_hd__buf_1 _11969_ (.A(_05951_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_2 _11970_ (.A0(_05744_),
    .A1(net576),
    .S(_05949_),
    .X(_05952_));
 sky130_fd_sc_hd__buf_1 _11971_ (.A(_05952_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_2 _11972_ (.A0(_04795_),
    .A1(net680),
    .S(_05949_),
    .X(_05953_));
 sky130_fd_sc_hd__buf_1 _11973_ (.A(_05953_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_2 _11974_ (.A0(_04801_),
    .A1(\rvsingle.dp.rf.rf[4][13] ),
    .S(_05949_),
    .X(_05954_));
 sky130_fd_sc_hd__buf_1 _11975_ (.A(_05954_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_2 _11976_ (.A0(_04807_),
    .A1(net400),
    .S(_05949_),
    .X(_05955_));
 sky130_fd_sc_hd__buf_1 _11977_ (.A(_05955_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_2 _11978_ (.A0(_04813_),
    .A1(net655),
    .S(_05949_),
    .X(_05956_));
 sky130_fd_sc_hd__buf_1 _11979_ (.A(_05956_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_2 _11980_ (.A0(_05344_),
    .A1(net386),
    .S(_05949_),
    .X(_05957_));
 sky130_fd_sc_hd__buf_1 _11981_ (.A(_05957_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_2 _11982_ (.A0(_04823_),
    .A1(net321),
    .S(_05949_),
    .X(_05958_));
 sky130_fd_sc_hd__buf_1 _11983_ (.A(_05958_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_2 _11984_ (.A0(_05173_),
    .A1(net327),
    .S(_05949_),
    .X(_05959_));
 sky130_fd_sc_hd__buf_1 _11985_ (.A(_05959_),
    .X(_00673_));
 sky130_fd_sc_hd__buf_1 _11986_ (.A(_05939_),
    .X(_05960_));
 sky130_fd_sc_hd__mux2_2 _11987_ (.A0(_04833_),
    .A1(net241),
    .S(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__buf_1 _11988_ (.A(_05961_),
    .X(_00674_));
 sky130_fd_sc_hd__o2bb2ai_2 _11989_ (.A1_N(net182),
    .A2_N(_05940_),
    .B1(_05835_),
    .B2(_05513_),
    .Y(_00675_));
 sky130_fd_sc_hd__mux2_2 _11990_ (.A0(_04845_),
    .A1(net278),
    .S(_05960_),
    .X(_05962_));
 sky130_fd_sc_hd__buf_1 _11991_ (.A(_05962_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_2 _11992_ (.A0(_04852_),
    .A1(net354),
    .S(_05960_),
    .X(_05963_));
 sky130_fd_sc_hd__buf_1 _11993_ (.A(_05963_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_2 _11994_ (.A0(_05757_),
    .A1(\rvsingle.dp.rf.rf[4][23] ),
    .S(_05960_),
    .X(_05964_));
 sky130_fd_sc_hd__buf_1 _11995_ (.A(_05964_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_2 _11996_ (.A0(_05132_),
    .A1(net375),
    .S(_05960_),
    .X(_05965_));
 sky130_fd_sc_hd__buf_1 _11997_ (.A(_05965_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_2 _11998_ (.A0(_04869_),
    .A1(net293),
    .S(_05960_),
    .X(_05966_));
 sky130_fd_sc_hd__buf_1 _11999_ (.A(_05966_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_2 _12000_ (.A0(_04876_),
    .A1(net262),
    .S(_05960_),
    .X(_05967_));
 sky130_fd_sc_hd__buf_1 _12001_ (.A(_05967_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_2 _12002_ (.A0(_05713_),
    .A1(net225),
    .S(_05960_),
    .X(_05968_));
 sky130_fd_sc_hd__buf_1 _12003_ (.A(_05968_),
    .X(_00682_));
 sky130_fd_sc_hd__a2bb2o_2 _12004_ (.A1_N(_05137_),
    .A2_N(_05847_),
    .B1(_05940_),
    .B2(net252),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_2 _12005_ (.A0(_05716_),
    .A1(net239),
    .S(_05960_),
    .X(_05969_));
 sky130_fd_sc_hd__buf_1 _12006_ (.A(_05969_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_2 _12007_ (.A0(_05639_),
    .A1(net243),
    .S(_05960_),
    .X(_05970_));
 sky130_fd_sc_hd__buf_1 _12008_ (.A(_05970_),
    .X(_00685_));
 sky130_fd_sc_hd__inv_2 _12009_ (.A(net29),
    .Y(_05971_));
 sky130_fd_sc_hd__o21ai_2 _12010_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05937_),
    .Y(_05972_));
 sky130_fd_sc_hd__o21ai_2 _12011_ (.A1(_05971_),
    .A2(_05937_),
    .B1(_05972_),
    .Y(_00686_));
 sky130_fd_sc_hd__and3_2 _12012_ (.A(_04721_),
    .B(_04920_),
    .C(_05142_),
    .X(_05973_));
 sky130_fd_sc_hd__a21oi_2 _12013_ (.A1(_05099_),
    .A2(_05146_),
    .B1(net149),
    .Y(_05974_));
 sky130_fd_sc_hd__a21oi_2 _12014_ (.A1(_05721_),
    .A2(_05973_),
    .B1(_05974_),
    .Y(_00687_));
 sky130_fd_sc_hd__or4_2 _12015_ (.A(_04737_),
    .B(_04919_),
    .C(_04733_),
    .D(_05149_),
    .X(_05975_));
 sky130_fd_sc_hd__buf_1 _12016_ (.A(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__mux2_2 _12017_ (.A0(_05724_),
    .A1(net578),
    .S(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__buf_1 _12018_ (.A(_05977_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_2 _12019_ (.A0(_05728_),
    .A1(net607),
    .S(_05976_),
    .X(_05978_));
 sky130_fd_sc_hd__buf_1 _12020_ (.A(_05978_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_2 _12021_ (.A0(_05531_),
    .A1(\rvsingle.dp.rf.rf[8][3] ),
    .S(_05976_),
    .X(_05979_));
 sky130_fd_sc_hd__buf_1 _12022_ (.A(_05979_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_2 _12023_ (.A0(_04759_),
    .A1(net396),
    .S(_05976_),
    .X(_05980_));
 sky130_fd_sc_hd__buf_1 _12024_ (.A(_05980_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_2 _12025_ (.A0(_04764_),
    .A1(net585),
    .S(_05976_),
    .X(_05981_));
 sky130_fd_sc_hd__buf_1 _12026_ (.A(_05981_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_2 _12027_ (.A0(_04769_),
    .A1(net390),
    .S(_05976_),
    .X(_05982_));
 sky130_fd_sc_hd__buf_1 _12028_ (.A(_05982_),
    .X(_00693_));
 sky130_fd_sc_hd__buf_1 _12029_ (.A(_05975_),
    .X(_05983_));
 sky130_fd_sc_hd__mux2_2 _12030_ (.A0(_04773_),
    .A1(net792),
    .S(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__buf_1 _12031_ (.A(_05984_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_2 _12032_ (.A0(_05740_),
    .A1(net777),
    .S(_05983_),
    .X(_05985_));
 sky130_fd_sc_hd__buf_1 _12033_ (.A(_05985_),
    .X(_00695_));
 sky130_fd_sc_hd__a22o_2 _12034_ (.A1(_05976_),
    .A2(net152),
    .B1(_05116_),
    .B2(_05146_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_2 _12035_ (.A0(_04785_),
    .A1(net613),
    .S(_05983_),
    .X(_05986_));
 sky130_fd_sc_hd__buf_1 _12036_ (.A(_05986_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_2 _12037_ (.A0(_05744_),
    .A1(net218),
    .S(_05983_),
    .X(_05987_));
 sky130_fd_sc_hd__buf_1 _12038_ (.A(_05987_),
    .X(_00698_));
 sky130_fd_sc_hd__a22o_2 _12039_ (.A1(_05976_),
    .A2(net168),
    .B1(_05119_),
    .B2(_05146_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_2 _12040_ (.A0(_04801_),
    .A1(net677),
    .S(_05983_),
    .X(_05988_));
 sky130_fd_sc_hd__buf_1 _12041_ (.A(_05988_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_2 _12042_ (.A0(_04807_),
    .A1(net530),
    .S(_05983_),
    .X(_05989_));
 sky130_fd_sc_hd__buf_1 _12043_ (.A(_05989_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_2 _12044_ (.A0(_04813_),
    .A1(net381),
    .S(_05983_),
    .X(_05990_));
 sky130_fd_sc_hd__buf_1 _12045_ (.A(_05990_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_2 _12046_ (.A0(_05344_),
    .A1(net537),
    .S(_05983_),
    .X(_05991_));
 sky130_fd_sc_hd__buf_1 _12047_ (.A(_05991_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_2 _12048_ (.A0(_04823_),
    .A1(net357),
    .S(_05983_),
    .X(_05992_));
 sky130_fd_sc_hd__buf_1 _12049_ (.A(_05992_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_2 _12050_ (.A0(_05173_),
    .A1(net476),
    .S(_05983_),
    .X(_05993_));
 sky130_fd_sc_hd__buf_1 _12051_ (.A(_05993_),
    .X(_00705_));
 sky130_fd_sc_hd__buf_1 _12052_ (.A(_05975_),
    .X(_05994_));
 sky130_fd_sc_hd__mux2_2 _12053_ (.A0(_04833_),
    .A1(net470),
    .S(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__buf_1 _12054_ (.A(_05995_),
    .X(_00706_));
 sky130_fd_sc_hd__o2bb2ai_2 _12055_ (.A1_N(_05976_),
    .A2_N(net161),
    .B1(_05149_),
    .B2(_05513_),
    .Y(_00707_));
 sky130_fd_sc_hd__mux2_2 _12056_ (.A0(_04845_),
    .A1(net666),
    .S(_05994_),
    .X(_05996_));
 sky130_fd_sc_hd__buf_1 _12057_ (.A(_05996_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_2 _12058_ (.A0(_04852_),
    .A1(net527),
    .S(_05994_),
    .X(_05997_));
 sky130_fd_sc_hd__buf_1 _12059_ (.A(_05997_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_2 _12060_ (.A0(_05757_),
    .A1(net242),
    .S(_05994_),
    .X(_05998_));
 sky130_fd_sc_hd__buf_1 _12061_ (.A(_05998_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_2 _12062_ (.A0(_05132_),
    .A1(net409),
    .S(_05994_),
    .X(_05999_));
 sky130_fd_sc_hd__buf_1 _12063_ (.A(_05999_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_2 _12064_ (.A0(_04869_),
    .A1(net727),
    .S(_05994_),
    .X(_06000_));
 sky130_fd_sc_hd__buf_1 _12065_ (.A(_06000_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_2 _12066_ (.A0(_04876_),
    .A1(net466),
    .S(_05994_),
    .X(_06001_));
 sky130_fd_sc_hd__buf_1 _12067_ (.A(_06001_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_2 _12068_ (.A0(_05713_),
    .A1(net814),
    .S(_05994_),
    .X(_06002_));
 sky130_fd_sc_hd__buf_1 _12069_ (.A(_06002_),
    .X(_00714_));
 sky130_fd_sc_hd__a2bb2o_2 _12070_ (.A1_N(_05137_),
    .A2_N(_05167_),
    .B1(_05976_),
    .B2(net358),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_2 _12071_ (.A0(_05716_),
    .A1(net288),
    .S(_05994_),
    .X(_06003_));
 sky130_fd_sc_hd__buf_1 _12072_ (.A(_06003_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_2 _12073_ (.A0(_05639_),
    .A1(net247),
    .S(_05994_),
    .X(_06004_));
 sky130_fd_sc_hd__buf_1 _12074_ (.A(_06004_),
    .X(_00717_));
 sky130_fd_sc_hd__inv_2 _12075_ (.A(net49),
    .Y(_06005_));
 sky130_fd_sc_hd__o21ai_2 _12076_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05973_),
    .Y(_06006_));
 sky130_fd_sc_hd__o21ai_2 _12077_ (.A1(_06005_),
    .A2(_05973_),
    .B1(_06006_),
    .Y(_00718_));
 sky130_fd_sc_hd__and3_2 _12078_ (.A(_04721_),
    .B(_04726_),
    .C(_04924_),
    .X(_06007_));
 sky130_fd_sc_hd__a21oi_2 _12079_ (.A1(_05316_),
    .A2(_05099_),
    .B1(net147),
    .Y(_06008_));
 sky130_fd_sc_hd__a21oi_2 _12080_ (.A1(_05721_),
    .A2(_06007_),
    .B1(_06008_),
    .Y(_00719_));
 sky130_fd_sc_hd__or4b_2 _12081_ (.A(_04737_),
    .B(_04919_),
    .C(_04733_),
    .D_N(_04725_),
    .X(_06009_));
 sky130_fd_sc_hd__buf_1 _12082_ (.A(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__mux2_2 _12083_ (.A0(_05724_),
    .A1(net540),
    .S(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__buf_1 _12084_ (.A(_06011_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_2 _12085_ (.A0(_05728_),
    .A1(\rvsingle.dp.rf.rf[0][2] ),
    .S(_06010_),
    .X(_06012_));
 sky130_fd_sc_hd__buf_1 _12086_ (.A(_06012_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_2 _12087_ (.A0(_04754_),
    .A1(\rvsingle.dp.rf.rf[0][3] ),
    .S(_06010_),
    .X(_06013_));
 sky130_fd_sc_hd__buf_1 _12088_ (.A(_06013_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_2 _12089_ (.A0(_04759_),
    .A1(net629),
    .S(_06010_),
    .X(_06014_));
 sky130_fd_sc_hd__buf_1 _12090_ (.A(_06014_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_2 _12091_ (.A0(_04764_),
    .A1(\rvsingle.dp.rf.rf[0][5] ),
    .S(_06010_),
    .X(_06015_));
 sky130_fd_sc_hd__buf_1 _12092_ (.A(_06015_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_2 _12093_ (.A0(_04769_),
    .A1(\rvsingle.dp.rf.rf[0][6] ),
    .S(_06010_),
    .X(_06016_));
 sky130_fd_sc_hd__buf_1 _12094_ (.A(_06016_),
    .X(_00725_));
 sky130_fd_sc_hd__and2_2 _12095_ (.A(_04773_),
    .B(_04726_),
    .X(_06017_));
 sky130_fd_sc_hd__a32o_2 _12096_ (.A1(_06017_),
    .A2(_05060_),
    .A3(_04924_),
    .B1(_06010_),
    .B2(net33),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_2 _12097_ (.A0(_05740_),
    .A1(net356),
    .S(_06010_),
    .X(_06018_));
 sky130_fd_sc_hd__buf_1 _12098_ (.A(_06018_),
    .X(_00727_));
 sky130_fd_sc_hd__buf_1 _12099_ (.A(_06009_),
    .X(_06019_));
 sky130_fd_sc_hd__mux2_2 _12100_ (.A0(_04781_),
    .A1(net551),
    .S(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__buf_1 _12101_ (.A(_06020_),
    .X(_00728_));
 sky130_fd_sc_hd__and2_2 _12102_ (.A(_04785_),
    .B(_04726_),
    .X(_06021_));
 sky130_fd_sc_hd__a32o_2 _12103_ (.A1(_06021_),
    .A2(_05060_),
    .A3(_04924_),
    .B1(_06010_),
    .B2(net15),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_2 _12104_ (.A0(_05744_),
    .A1(net450),
    .S(_06019_),
    .X(_06022_));
 sky130_fd_sc_hd__buf_1 _12105_ (.A(_06022_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_2 _12106_ (.A0(_04795_),
    .A1(net513),
    .S(_06019_),
    .X(_06023_));
 sky130_fd_sc_hd__buf_1 _12107_ (.A(_06023_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_2 _12108_ (.A0(_04801_),
    .A1(net554),
    .S(_06019_),
    .X(_06024_));
 sky130_fd_sc_hd__buf_1 _12109_ (.A(_06024_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_2 _12110_ (.A0(_04807_),
    .A1(net531),
    .S(_06019_),
    .X(_06025_));
 sky130_fd_sc_hd__buf_1 _12111_ (.A(_06025_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_2 _12112_ (.A0(_04813_),
    .A1(net532),
    .S(_06019_),
    .X(_06026_));
 sky130_fd_sc_hd__buf_1 _12113_ (.A(_06026_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_2 _12114_ (.A0(_05344_),
    .A1(net428),
    .S(_06019_),
    .X(_06027_));
 sky130_fd_sc_hd__buf_1 _12115_ (.A(_06027_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_2 _12116_ (.A0(_04823_),
    .A1(net265),
    .S(_06019_),
    .X(_06028_));
 sky130_fd_sc_hd__buf_1 _12117_ (.A(_06028_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_2 _12118_ (.A0(_05173_),
    .A1(net642),
    .S(_06019_),
    .X(_06029_));
 sky130_fd_sc_hd__buf_1 _12119_ (.A(_06029_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_2 _12120_ (.A0(_04833_),
    .A1(net472),
    .S(_06019_),
    .X(_06030_));
 sky130_fd_sc_hd__buf_1 _12121_ (.A(_06030_),
    .X(_00738_));
 sky130_fd_sc_hd__buf_1 _12122_ (.A(_06009_),
    .X(_06031_));
 sky130_fd_sc_hd__mux2_2 _12123_ (.A0(_04839_),
    .A1(net674),
    .S(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__buf_1 _12124_ (.A(_06032_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_2 _12125_ (.A0(_04845_),
    .A1(net791),
    .S(_06031_),
    .X(_06033_));
 sky130_fd_sc_hd__buf_1 _12126_ (.A(_06033_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_2 _12127_ (.A0(_04852_),
    .A1(net398),
    .S(_06031_),
    .X(_06034_));
 sky130_fd_sc_hd__buf_1 _12128_ (.A(_06034_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_2 _12129_ (.A0(_05757_),
    .A1(net608),
    .S(_06031_),
    .X(_06035_));
 sky130_fd_sc_hd__buf_1 _12130_ (.A(_06035_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_2 _12131_ (.A0(_05132_),
    .A1(net348),
    .S(_06031_),
    .X(_06036_));
 sky130_fd_sc_hd__buf_1 _12132_ (.A(_06036_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_2 _12133_ (.A0(_04869_),
    .A1(net482),
    .S(_06031_),
    .X(_06037_));
 sky130_fd_sc_hd__buf_1 _12134_ (.A(_06037_),
    .X(_00744_));
 sky130_fd_sc_hd__and2_2 _12135_ (.A(_04876_),
    .B(_04726_),
    .X(_06038_));
 sky130_fd_sc_hd__a32o_2 _12136_ (.A1(_06038_),
    .A2(_05060_),
    .A3(_04924_),
    .B1(_06010_),
    .B2(net180),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_2 _12137_ (.A0(_05713_),
    .A1(net362),
    .S(_06031_),
    .X(_06039_));
 sky130_fd_sc_hd__buf_1 _12138_ (.A(_06039_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_2 _12139_ (.A0(_05763_),
    .A1(net331),
    .S(_06031_),
    .X(_06040_));
 sky130_fd_sc_hd__buf_1 _12140_ (.A(_06040_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_2 _12141_ (.A0(_05716_),
    .A1(net219),
    .S(_06031_),
    .X(_06041_));
 sky130_fd_sc_hd__buf_1 _12142_ (.A(_06041_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_2 _12143_ (.A0(_05639_),
    .A1(net267),
    .S(_06031_),
    .X(_06042_));
 sky130_fd_sc_hd__buf_1 _12144_ (.A(_06042_),
    .X(_00749_));
 sky130_fd_sc_hd__inv_2 _12145_ (.A(net61),
    .Y(_06043_));
 sky130_fd_sc_hd__o21ai_2 _12146_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_06007_),
    .Y(_06044_));
 sky130_fd_sc_hd__o21ai_2 _12147_ (.A1(_06043_),
    .A2(_06007_),
    .B1(_06044_),
    .Y(_00750_));
 sky130_fd_sc_hd__and4_2 _12148_ (.A(_04720_),
    .B(_04725_),
    .C(_04967_),
    .D(_04968_),
    .X(_06045_));
 sky130_fd_sc_hd__a21oi_2 _12149_ (.A1(_05316_),
    .A2(_04973_),
    .B1(net28),
    .Y(_06046_));
 sky130_fd_sc_hd__a21oi_2 _12150_ (.A1(_05721_),
    .A2(_06045_),
    .B1(_06046_),
    .Y(_00751_));
 sky130_fd_sc_hd__or4_2 _12151_ (.A(_04722_),
    .B(_04723_),
    .C(_04724_),
    .D(_05003_),
    .X(_06047_));
 sky130_fd_sc_hd__buf_1 _12152_ (.A(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__buf_1 _12153_ (.A(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__mux2_2 _12154_ (.A0(_05724_),
    .A1(net684),
    .S(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__buf_1 _12155_ (.A(_06050_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_2 _12156_ (.A0(_05728_),
    .A1(net775),
    .S(_06049_),
    .X(_06051_));
 sky130_fd_sc_hd__buf_1 _12157_ (.A(_06051_),
    .X(_00753_));
 sky130_fd_sc_hd__buf_1 _12158_ (.A(_06049_),
    .X(_06052_));
 sky130_fd_sc_hd__a2bb2o_2 _12159_ (.A1_N(_05004_),
    .A2_N(_05324_),
    .B1(_06052_),
    .B2(net138),
    .X(_00754_));
 sky130_fd_sc_hd__a2bb2o_2 _12160_ (.A1_N(_05004_),
    .A2_N(_05326_),
    .B1(_06052_),
    .B2(net203),
    .X(_00755_));
 sky130_fd_sc_hd__a22o_2 _12161_ (.A1(net100),
    .A2(_06052_),
    .B1(_05327_),
    .B2(_04985_),
    .X(_00756_));
 sky130_fd_sc_hd__a2bb2o_2 _12162_ (.A1_N(_05004_),
    .A2_N(_05328_),
    .B1(_06052_),
    .B2(net211),
    .X(_00757_));
 sky130_fd_sc_hd__a22o_2 _12163_ (.A1(net19),
    .A2(_06052_),
    .B1(_06017_),
    .B2(_04985_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_2 _12164_ (.A0(_05740_),
    .A1(net511),
    .S(_06049_),
    .X(_06053_));
 sky130_fd_sc_hd__buf_1 _12165_ (.A(_06053_),
    .X(_00759_));
 sky130_fd_sc_hd__a22o_2 _12166_ (.A1(net21),
    .A2(_06052_),
    .B1(_05332_),
    .B2(_04985_),
    .X(_00760_));
 sky130_fd_sc_hd__a22o_2 _12167_ (.A1(net85),
    .A2(_06049_),
    .B1(_06021_),
    .B2(_04985_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_2 _12168_ (.A0(_05744_),
    .A1(net224),
    .S(_06049_),
    .X(_06054_));
 sky130_fd_sc_hd__buf_1 _12169_ (.A(_06054_),
    .X(_00762_));
 sky130_fd_sc_hd__o41a_2 _12170_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05004_),
    .B1(net194),
    .X(_06055_));
 sky130_fd_sc_hd__a31o_2 _12171_ (.A1(_04796_),
    .A2(_05766_),
    .A3(_05336_),
    .B1(_06055_),
    .X(_00763_));
 sky130_fd_sc_hd__o41a_2 _12172_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05003_),
    .B1(net201),
    .X(_06056_));
 sky130_fd_sc_hd__a31o_2 _12173_ (.A1(_04802_),
    .A2(_05766_),
    .A3(_05336_),
    .B1(_06056_),
    .X(_00764_));
 sky130_fd_sc_hd__a2bb2o_2 _12174_ (.A1_N(_05004_),
    .A2_N(_05342_),
    .B1(_06052_),
    .B2(net97),
    .X(_00765_));
 sky130_fd_sc_hd__a2bb2o_2 _12175_ (.A1_N(_05004_),
    .A2_N(_05343_),
    .B1(_06052_),
    .B2(net151),
    .X(_00766_));
 sky130_fd_sc_hd__a22o_2 _12176_ (.A1(net176),
    .A2(_06049_),
    .B1(_05345_),
    .B2(_04985_),
    .X(_00767_));
 sky130_fd_sc_hd__a22o_2 _12177_ (.A1(net103),
    .A2(_06049_),
    .B1(_05346_),
    .B2(_05766_),
    .X(_00768_));
 sky130_fd_sc_hd__a22o_2 _12178_ (.A1(net20),
    .A2(_06049_),
    .B1(_05347_),
    .B2(_05766_),
    .X(_00769_));
 sky130_fd_sc_hd__a2bb2o_2 _12179_ (.A1_N(_05004_),
    .A2_N(_05348_),
    .B1(_06052_),
    .B2(net174),
    .X(_00770_));
 sky130_fd_sc_hd__o41a_2 _12180_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05003_),
    .B1(net192),
    .X(_06057_));
 sky130_fd_sc_hd__a31o_2 _12181_ (.A1(_04840_),
    .A2(_05766_),
    .A3(_05336_),
    .B1(_06057_),
    .X(_00771_));
 sky130_fd_sc_hd__a2bb2o_2 _12182_ (.A1_N(_05004_),
    .A2_N(_05350_),
    .B1(_06052_),
    .B2(net177),
    .X(_00772_));
 sky130_fd_sc_hd__o41a_2 _12183_ (.A1(_05337_),
    .A2(_05338_),
    .A3(_05339_),
    .A4(_05003_),
    .B1(net207),
    .X(_06058_));
 sky130_fd_sc_hd__a31o_2 _12184_ (.A1(_04853_),
    .A2(_05766_),
    .A3(_05336_),
    .B1(_06058_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_2 _12185_ (.A0(_05757_),
    .A1(net307),
    .S(_06048_),
    .X(_06059_));
 sky130_fd_sc_hd__buf_1 _12186_ (.A(_06059_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_2 _12187_ (.A0(_05132_),
    .A1(net378),
    .S(_06048_),
    .X(_06060_));
 sky130_fd_sc_hd__buf_1 _12188_ (.A(_06060_),
    .X(_00775_));
 sky130_fd_sc_hd__o41a_2 _12189_ (.A1(_04982_),
    .A2(_04983_),
    .A3(_04981_),
    .A4(_05003_),
    .B1(net388),
    .X(_06061_));
 sky130_fd_sc_hd__a31o_2 _12190_ (.A1(_04870_),
    .A2(_05766_),
    .A3(_05316_),
    .B1(_06061_),
    .X(_00776_));
 sky130_fd_sc_hd__a22o_2 _12191_ (.A1(net141),
    .A2(_06049_),
    .B1(_06038_),
    .B2(_05766_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_2 _12192_ (.A0(_04885_),
    .A1(\rvsingle.dp.rf.rf[3][27] ),
    .S(_06048_),
    .X(_06062_));
 sky130_fd_sc_hd__buf_1 _12193_ (.A(_06062_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_2 _12194_ (.A0(_05763_),
    .A1(net324),
    .S(_06048_),
    .X(_06063_));
 sky130_fd_sc_hd__buf_1 _12195_ (.A(_06063_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_2 _12196_ (.A0(_04897_),
    .A1(net667),
    .S(_06048_),
    .X(_06064_));
 sky130_fd_sc_hd__buf_1 _12197_ (.A(_06064_),
    .X(_00780_));
 sky130_fd_sc_hd__o41a_2 _12198_ (.A1(_04982_),
    .A2(_04983_),
    .A3(_04981_),
    .A4(_05003_),
    .B1(net313),
    .X(_06065_));
 sky130_fd_sc_hd__a31o_2 _12199_ (.A1(_04904_),
    .A2(_04973_),
    .A3(_05316_),
    .B1(_06065_),
    .X(_00781_));
 sky130_fd_sc_hd__inv_2 _12200_ (.A(net62),
    .Y(_06066_));
 sky130_fd_sc_hd__o21ai_2 _12201_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_06045_),
    .Y(_06067_));
 sky130_fd_sc_hd__o21ai_2 _12202_ (.A1(_06066_),
    .A2(_06045_),
    .B1(_06067_),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _12203_ (.A(_05898_),
    .Y(_00002_));
 sky130_fd_sc_hd__inv_2 _12204_ (.A(_05898_),
    .Y(_00003_));
 sky130_fd_sc_hd__inv_2 _12205_ (.A(_05898_),
    .Y(_00004_));
 sky130_fd_sc_hd__inv_2 _12206_ (.A(_05898_),
    .Y(_00005_));
 sky130_fd_sc_hd__inv_2 _12207_ (.A(_05898_),
    .Y(_00006_));
 sky130_fd_sc_hd__inv_2 _12208_ (.A(_05898_),
    .Y(_00007_));
 sky130_fd_sc_hd__inv_2 _12209_ (.A(_05898_),
    .Y(_00008_));
 sky130_fd_sc_hd__inv_2 _12210_ (.A(_05898_),
    .Y(_00009_));
 sky130_fd_sc_hd__buf_1 _12211_ (.A(reset),
    .X(_06068_));
 sky130_fd_sc_hd__inv_2 _12212_ (.A(_06068_),
    .Y(_00010_));
 sky130_fd_sc_hd__inv_2 _12213_ (.A(_06068_),
    .Y(_00011_));
 sky130_fd_sc_hd__inv_2 _12214_ (.A(_06068_),
    .Y(_00012_));
 sky130_fd_sc_hd__inv_2 _12215_ (.A(_06068_),
    .Y(_00013_));
 sky130_fd_sc_hd__inv_2 _12216_ (.A(_06068_),
    .Y(_00014_));
 sky130_fd_sc_hd__inv_2 _12217_ (.A(_06068_),
    .Y(_00015_));
 sky130_fd_sc_hd__inv_2 _12218_ (.A(_06068_),
    .Y(_00016_));
 sky130_fd_sc_hd__inv_2 _12219_ (.A(_06068_),
    .Y(_00017_));
 sky130_fd_sc_hd__inv_2 _12220_ (.A(_06068_),
    .Y(_00018_));
 sky130_fd_sc_hd__inv_2 _12221_ (.A(_06068_),
    .Y(_00019_));
 sky130_fd_sc_hd__buf_1 _12222_ (.A(reset),
    .X(_06069_));
 sky130_fd_sc_hd__inv_2 _12223_ (.A(_06069_),
    .Y(_00020_));
 sky130_fd_sc_hd__inv_2 _12224_ (.A(_06069_),
    .Y(_00021_));
 sky130_fd_sc_hd__inv_2 _12225_ (.A(_06069_),
    .Y(_00022_));
 sky130_fd_sc_hd__inv_2 _12226_ (.A(_06069_),
    .Y(_00023_));
 sky130_fd_sc_hd__inv_2 _12227_ (.A(_06069_),
    .Y(_00024_));
 sky130_fd_sc_hd__inv_2 _12228_ (.A(_06069_),
    .Y(_00025_));
 sky130_fd_sc_hd__inv_2 _12229_ (.A(_06069_),
    .Y(_00026_));
 sky130_fd_sc_hd__inv_2 _12230_ (.A(_06069_),
    .Y(_00027_));
 sky130_fd_sc_hd__inv_2 _12231_ (.A(_06069_),
    .Y(_00028_));
 sky130_fd_sc_hd__inv_2 _12232_ (.A(_06069_),
    .Y(_00029_));
 sky130_fd_sc_hd__inv_2 _12233_ (.A(reset),
    .Y(_00030_));
 sky130_fd_sc_hd__inv_2 _12234_ (.A(reset),
    .Y(_00031_));
 sky130_fd_sc_hd__and3_2 _12235_ (.A(_04721_),
    .B(_05058_),
    .C(_05830_),
    .X(_06070_));
 sky130_fd_sc_hd__a21oi_2 _12236_ (.A1(_05145_),
    .A2(_05830_),
    .B1(net164),
    .Y(_06071_));
 sky130_fd_sc_hd__a21oi_2 _12237_ (.A1(_04718_),
    .A2(_06070_),
    .B1(_06071_),
    .Y(_00783_));
 sky130_fd_sc_hd__or4b_2 _12238_ (.A(_04919_),
    .B(_04732_),
    .C(_05835_),
    .D_N(_04737_),
    .X(_06072_));
 sky130_fd_sc_hd__buf_1 _12239_ (.A(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__buf_1 _12240_ (.A(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__mux2_2 _12241_ (.A0(_04735_),
    .A1(\rvsingle.dp.rf.rf[5][1] ),
    .S(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__buf_1 _12242_ (.A(_06075_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_2 _12243_ (.A0(_04746_),
    .A1(net636),
    .S(_06074_),
    .X(_06076_));
 sky130_fd_sc_hd__buf_1 _12244_ (.A(_06076_),
    .X(_00785_));
 sky130_fd_sc_hd__buf_1 _12245_ (.A(_06074_),
    .X(_06077_));
 sky130_fd_sc_hd__a22o_2 _12246_ (.A1(_06077_),
    .A2(net45),
    .B1(_05156_),
    .B2(_05841_),
    .X(_00786_));
 sky130_fd_sc_hd__a22o_2 _12247_ (.A1(_06077_),
    .A2(net181),
    .B1(_05465_),
    .B2(_05832_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_2 _12248_ (.A0(_04764_),
    .A1(\rvsingle.dp.rf.rf[5][5] ),
    .S(_06074_),
    .X(_06078_));
 sky130_fd_sc_hd__buf_1 _12249_ (.A(_06078_),
    .X(_00788_));
 sky130_fd_sc_hd__a22o_2 _12250_ (.A1(_06077_),
    .A2(net129),
    .B1(_05466_),
    .B2(_05832_),
    .X(_00789_));
 sky130_fd_sc_hd__a22o_2 _12251_ (.A1(_06077_),
    .A2(net89),
    .B1(_05161_),
    .B2(_05832_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_2 _12252_ (.A0(_04777_),
    .A1(\rvsingle.dp.rf.rf[5][8] ),
    .S(_06074_),
    .X(_06079_));
 sky130_fd_sc_hd__buf_1 _12253_ (.A(_06079_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_2 _12254_ (.A0(_04781_),
    .A1(\rvsingle.dp.rf.rf[5][9] ),
    .S(_06074_),
    .X(_06080_));
 sky130_fd_sc_hd__buf_1 _12255_ (.A(_06080_),
    .X(_00792_));
 sky130_fd_sc_hd__a22o_2 _12256_ (.A1(_06077_),
    .A2(net52),
    .B1(_05164_),
    .B2(_05832_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_2 _12257_ (.A0(_05744_),
    .A1(net231),
    .S(_06074_),
    .X(_06081_));
 sky130_fd_sc_hd__buf_1 _12258_ (.A(_06081_),
    .X(_00794_));
 sky130_fd_sc_hd__a2bb2o_2 _12259_ (.A1_N(_05472_),
    .A2_N(_05847_),
    .B1(_06077_),
    .B2(net170),
    .X(_00795_));
 sky130_fd_sc_hd__a2bb2o_2 _12260_ (.A1_N(_05168_),
    .A2_N(_05847_),
    .B1(_06077_),
    .B2(net128),
    .X(_00796_));
 sky130_fd_sc_hd__a2bb2o_2 _12261_ (.A1_N(_05169_),
    .A2_N(_05847_),
    .B1(_06077_),
    .B2(net83),
    .X(_00797_));
 sky130_fd_sc_hd__a2bb2o_2 _12262_ (.A1_N(_05474_),
    .A2_N(_05847_),
    .B1(_06077_),
    .B2(net82),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_2 _12263_ (.A0(_05344_),
    .A1(net232),
    .S(_06074_),
    .X(_06082_));
 sky130_fd_sc_hd__buf_1 _12264_ (.A(_06082_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_2 _12265_ (.A0(_04823_),
    .A1(net435),
    .S(_06073_),
    .X(_06083_));
 sky130_fd_sc_hd__buf_1 _12266_ (.A(_06083_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_2 _12267_ (.A0(_05173_),
    .A1(net494),
    .S(_06073_),
    .X(_06084_));
 sky130_fd_sc_hd__buf_1 _12268_ (.A(_06084_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_2 _12269_ (.A0(_04833_),
    .A1(net439),
    .S(_06073_),
    .X(_06085_));
 sky130_fd_sc_hd__buf_1 _12270_ (.A(_06085_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_2 _12271_ (.A0(_04839_),
    .A1(net316),
    .S(_06073_),
    .X(_06086_));
 sky130_fd_sc_hd__buf_1 _12272_ (.A(_06086_),
    .X(_00803_));
 sky130_fd_sc_hd__a2bb2o_2 _12273_ (.A1_N(_05177_),
    .A2_N(_05835_),
    .B1(_06077_),
    .B2(net171),
    .X(_00804_));
 sky130_fd_sc_hd__a22o_2 _12274_ (.A1(_06074_),
    .A2(net96),
    .B1(_05178_),
    .B2(_05832_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_2 _12275_ (.A0(_04858_),
    .A1(net596),
    .S(_06073_),
    .X(_06087_));
 sky130_fd_sc_hd__buf_1 _12276_ (.A(_06087_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_2 _12277_ (.A0(_05132_),
    .A1(net303),
    .S(_06073_),
    .X(_06088_));
 sky130_fd_sc_hd__buf_1 _12278_ (.A(_06088_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_2 _12279_ (.A0(_04869_),
    .A1(net620),
    .S(_06073_),
    .X(_06089_));
 sky130_fd_sc_hd__buf_1 _12280_ (.A(_06089_),
    .X(_00808_));
 sky130_fd_sc_hd__a22o_2 _12281_ (.A1(_06074_),
    .A2(net134),
    .B1(_05182_),
    .B2(_05832_),
    .X(_00809_));
 sky130_fd_sc_hd__o21a_2 _12282_ (.A1(_05084_),
    .A2(_05835_),
    .B1(net215),
    .X(_06090_));
 sky130_fd_sc_hd__a31o_2 _12283_ (.A1(_04886_),
    .A2(_05183_),
    .A3(_05832_),
    .B1(_06090_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_2 _12284_ (.A0(_05763_),
    .A1(net264),
    .S(_06073_),
    .X(_06091_));
 sky130_fd_sc_hd__buf_1 _12285_ (.A(_06091_),
    .X(_00811_));
 sky130_fd_sc_hd__o21a_2 _12286_ (.A1(_05084_),
    .A2(_05835_),
    .B1(net276),
    .X(_06092_));
 sky130_fd_sc_hd__a31o_2 _12287_ (.A1(_04898_),
    .A2(_05145_),
    .A3(_05832_),
    .B1(_06092_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_2 _12288_ (.A0(_04903_),
    .A1(net474),
    .S(_06073_),
    .X(_06093_));
 sky130_fd_sc_hd__buf_1 _12289_ (.A(_06093_),
    .X(_00813_));
 sky130_fd_sc_hd__inv_2 _12290_ (.A(net90),
    .Y(_06094_));
 sky130_fd_sc_hd__o21ai_2 _12291_ (.A1(_04908_),
    .A2(_04912_),
    .B1(_06070_),
    .Y(_06095_));
 sky130_fd_sc_hd__o21ai_2 _12292_ (.A1(_06094_),
    .A2(_06070_),
    .B1(_06095_),
    .Y(_00814_));
 sky130_fd_sc_hd__and4_2 _12293_ (.A(_04916_),
    .B(_04918_),
    .C(_04728_),
    .D(_04922_),
    .X(_06096_));
 sky130_fd_sc_hd__a21oi_2 _12294_ (.A1(_04728_),
    .A2(_04925_),
    .B1(net53),
    .Y(_06097_));
 sky130_fd_sc_hd__a21oi_2 _12295_ (.A1(_04718_),
    .A2(_06096_),
    .B1(_06097_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_2 _12296_ (.A(_04728_),
    .B(_04925_),
    .Y(_06098_));
 sky130_fd_sc_hd__buf_1 _12297_ (.A(_06098_),
    .X(_06099_));
 sky130_fd_sc_hd__mux2_2 _12298_ (.A0(_04735_),
    .A1(\rvsingle.dp.rf.rf[30][1] ),
    .S(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__buf_1 _12299_ (.A(_06100_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_2 _12300_ (.A0(_04746_),
    .A1(\rvsingle.dp.rf.rf[30][2] ),
    .S(_06099_),
    .X(_06101_));
 sky130_fd_sc_hd__buf_1 _12301_ (.A(_06101_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_2 _12302_ (.A0(_04754_),
    .A1(net610),
    .S(_06099_),
    .X(_06102_));
 sky130_fd_sc_hd__buf_1 _12303_ (.A(_06102_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_2 _12304_ (.A0(_04759_),
    .A1(net706),
    .S(_06099_),
    .X(_06103_));
 sky130_fd_sc_hd__buf_1 _12305_ (.A(_06103_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_2 _12306_ (.A0(_04764_),
    .A1(net481),
    .S(_06099_),
    .X(_06104_));
 sky130_fd_sc_hd__buf_1 _12307_ (.A(_06104_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_2 _12308_ (.A0(_04769_),
    .A1(net749),
    .S(_06099_),
    .X(_06105_));
 sky130_fd_sc_hd__buf_1 _12309_ (.A(_06105_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_2 _12310_ (.A0(_04773_),
    .A1(net622),
    .S(_06099_),
    .X(_06106_));
 sky130_fd_sc_hd__buf_1 _12311_ (.A(_06106_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_2 _12312_ (.A0(_04777_),
    .A1(\rvsingle.dp.rf.rf[30][8] ),
    .S(_06099_),
    .X(_06107_));
 sky130_fd_sc_hd__buf_1 _12313_ (.A(_06107_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_2 _12314_ (.A0(_04781_),
    .A1(net599),
    .S(_06099_),
    .X(_06108_));
 sky130_fd_sc_hd__buf_1 _12315_ (.A(_06108_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_2 _12316_ (.A0(_04785_),
    .A1(net525),
    .S(_06099_),
    .X(_06109_));
 sky130_fd_sc_hd__buf_1 _12317_ (.A(_06109_),
    .X(_00825_));
 sky130_fd_sc_hd__buf_1 _12318_ (.A(_06098_),
    .X(_06110_));
 sky130_fd_sc_hd__mux2_2 _12319_ (.A0(_05744_),
    .A1(net284),
    .S(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__buf_1 _12320_ (.A(_06111_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_2 _12321_ (.A0(_04795_),
    .A1(net506),
    .S(_06110_),
    .X(_06112_));
 sky130_fd_sc_hd__buf_1 _12322_ (.A(_06112_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_2 _12323_ (.A0(_04801_),
    .A1(net593),
    .S(_06110_),
    .X(_06113_));
 sky130_fd_sc_hd__buf_1 _12324_ (.A(_06113_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_2 _12325_ (.A0(_04807_),
    .A1(net804),
    .S(_06110_),
    .X(_06114_));
 sky130_fd_sc_hd__buf_1 _12326_ (.A(_06114_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_2 _12327_ (.A0(_04813_),
    .A1(net688),
    .S(_06110_),
    .X(_06115_));
 sky130_fd_sc_hd__buf_1 _12328_ (.A(_06115_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_2 _12329_ (.A0(_05344_),
    .A1(net490),
    .S(_06110_),
    .X(_06116_));
 sky130_fd_sc_hd__buf_1 _12330_ (.A(_06116_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_2 _12331_ (.A0(_04823_),
    .A1(net373),
    .S(_06110_),
    .X(_06117_));
 sky130_fd_sc_hd__buf_1 _12332_ (.A(_06117_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_2 _12333_ (.A0(_05173_),
    .A1(net760),
    .S(_06110_),
    .X(_06118_));
 sky130_fd_sc_hd__buf_1 _12334_ (.A(_06118_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_2 _12335_ (.A0(_04833_),
    .A1(net651),
    .S(_06110_),
    .X(_06119_));
 sky130_fd_sc_hd__buf_1 _12336_ (.A(_06119_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_2 _12337_ (.A0(_04839_),
    .A1(net700),
    .S(_06110_),
    .X(_06120_));
 sky130_fd_sc_hd__buf_1 _12338_ (.A(_06120_),
    .X(_00835_));
 sky130_fd_sc_hd__buf_1 _12339_ (.A(_06098_),
    .X(_06121_));
 sky130_fd_sc_hd__mux2_2 _12340_ (.A0(_04845_),
    .A1(net716),
    .S(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__buf_1 _12341_ (.A(_06122_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_2 _12342_ (.A0(_04852_),
    .A1(net574),
    .S(_06121_),
    .X(_06123_));
 sky130_fd_sc_hd__buf_1 _12343_ (.A(_06123_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_2 _12344_ (.A0(_04858_),
    .A1(net226),
    .S(_06121_),
    .X(_06124_));
 sky130_fd_sc_hd__buf_1 _12345_ (.A(_06124_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_2 _12346_ (.A0(_05132_),
    .A1(net401),
    .S(_06121_),
    .X(_06125_));
 sky130_fd_sc_hd__buf_1 _12347_ (.A(_06125_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_2 _12348_ (.A0(_04869_),
    .A1(net475),
    .S(_06121_),
    .X(_06126_));
 sky130_fd_sc_hd__buf_1 _12349_ (.A(_06126_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_2 _12350_ (.A0(_04876_),
    .A1(net268),
    .S(_06121_),
    .X(_06127_));
 sky130_fd_sc_hd__buf_1 _12351_ (.A(_06127_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_2 _12352_ (.A0(_04885_),
    .A1(net305),
    .S(_06121_),
    .X(_06128_));
 sky130_fd_sc_hd__buf_1 _12353_ (.A(_06128_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_2 _12354_ (.A0(_05763_),
    .A1(net221),
    .S(_06121_),
    .X(_06129_));
 sky130_fd_sc_hd__buf_1 _12355_ (.A(_06129_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_2 _12356_ (.A0(_04897_),
    .A1(net261),
    .S(_06121_),
    .X(_06130_));
 sky130_fd_sc_hd__buf_1 _12357_ (.A(_06130_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_2 _12358_ (.A0(_04903_),
    .A1(net258),
    .S(_06121_),
    .X(_06131_));
 sky130_fd_sc_hd__buf_1 _12359_ (.A(_06131_),
    .X(_00845_));
 sky130_fd_sc_hd__inv_2 _12360_ (.A(net25),
    .Y(_06132_));
 sky130_fd_sc_hd__o21ai_2 _12361_ (.A1(_04908_),
    .A2(_04912_),
    .B1(_06096_),
    .Y(_06133_));
 sky130_fd_sc_hd__o21ai_2 _12362_ (.A1(_06132_),
    .A2(_06096_),
    .B1(_06133_),
    .Y(_00846_));
 sky130_fd_sc_hd__dfxtp_2 _12363_ (.CLK(clknet_leaf_88_clk),
    .D(_00847_),
    .Q(\rvsingle.dp.rf.rf[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12364_ (.CLK(clknet_leaf_52_clk),
    .D(_00848_),
    .Q(\rvsingle.dp.rf.rf[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12365_ (.CLK(clknet_leaf_44_clk),
    .D(_00849_),
    .Q(\rvsingle.dp.rf.rf[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12366_ (.CLK(clknet_leaf_71_clk),
    .D(_00850_),
    .Q(\rvsingle.dp.rf.rf[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12367_ (.CLK(clknet_leaf_57_clk),
    .D(_00851_),
    .Q(\rvsingle.dp.rf.rf[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12368_ (.CLK(clknet_leaf_72_clk),
    .D(_00852_),
    .Q(\rvsingle.dp.rf.rf[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12369_ (.CLK(clknet_leaf_49_clk),
    .D(_00853_),
    .Q(\rvsingle.dp.rf.rf[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12370_ (.CLK(clknet_leaf_57_clk),
    .D(_00854_),
    .Q(\rvsingle.dp.rf.rf[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12371_ (.CLK(clknet_leaf_29_clk),
    .D(_00855_),
    .Q(\rvsingle.dp.rf.rf[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12372_ (.CLK(clknet_leaf_21_clk),
    .D(_00856_),
    .Q(\rvsingle.dp.rf.rf[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12373_ (.CLK(clknet_leaf_60_clk),
    .D(_00857_),
    .Q(\rvsingle.dp.rf.rf[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12374_ (.CLK(clknet_leaf_25_clk),
    .D(_00858_),
    .Q(\rvsingle.dp.rf.rf[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12375_ (.CLK(clknet_leaf_18_clk),
    .D(_00859_),
    .Q(\rvsingle.dp.rf.rf[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12376_ (.CLK(clknet_leaf_18_clk),
    .D(_00860_),
    .Q(\rvsingle.dp.rf.rf[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12377_ (.CLK(clknet_leaf_17_clk),
    .D(_00861_),
    .Q(\rvsingle.dp.rf.rf[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12378_ (.CLK(clknet_leaf_14_clk),
    .D(_00862_),
    .Q(\rvsingle.dp.rf.rf[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12379_ (.CLK(clknet_leaf_136_clk),
    .D(_00863_),
    .Q(\rvsingle.dp.rf.rf[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12380_ (.CLK(clknet_leaf_147_clk),
    .D(_00864_),
    .Q(\rvsingle.dp.rf.rf[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12381_ (.CLK(clknet_leaf_135_clk),
    .D(_00865_),
    .Q(\rvsingle.dp.rf.rf[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12382_ (.CLK(clknet_leaf_133_clk),
    .D(_00866_),
    .Q(\rvsingle.dp.rf.rf[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12383_ (.CLK(clknet_leaf_132_clk),
    .D(_00867_),
    .Q(\rvsingle.dp.rf.rf[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12384_ (.CLK(clknet_leaf_119_clk),
    .D(_00868_),
    .Q(\rvsingle.dp.rf.rf[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12385_ (.CLK(clknet_leaf_125_clk),
    .D(_00869_),
    .Q(\rvsingle.dp.rf.rf[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12386_ (.CLK(clknet_leaf_130_clk),
    .D(_00870_),
    .Q(\rvsingle.dp.rf.rf[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12387_ (.CLK(clknet_leaf_125_clk),
    .D(_00871_),
    .Q(\rvsingle.dp.rf.rf[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12388_ (.CLK(clknet_leaf_122_clk),
    .D(_00872_),
    .Q(\rvsingle.dp.rf.rf[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12389_ (.CLK(clknet_leaf_111_clk),
    .D(_00873_),
    .Q(\rvsingle.dp.rf.rf[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12390_ (.CLK(clknet_leaf_121_clk),
    .D(_00874_),
    .Q(\rvsingle.dp.rf.rf[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12391_ (.CLK(clknet_leaf_99_clk),
    .D(_00875_),
    .Q(\rvsingle.dp.rf.rf[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12392_ (.CLK(clknet_leaf_104_clk),
    .D(_00876_),
    .Q(\rvsingle.dp.rf.rf[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12393_ (.CLK(clknet_leaf_92_clk),
    .D(_00877_),
    .Q(\rvsingle.dp.rf.rf[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12394_ (.CLK(clknet_leaf_83_clk),
    .D(_00878_),
    .Q(\rvsingle.dp.rf.rf[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12395_ (.CLK(clknet_leaf_87_clk),
    .D(_00879_),
    .Q(\rvsingle.dp.rf.rf[28][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12396_ (.CLK(clknet_leaf_50_clk),
    .D(_00880_),
    .Q(\rvsingle.dp.rf.rf[28][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12397_ (.CLK(clknet_leaf_43_clk),
    .D(_00881_),
    .Q(\rvsingle.dp.rf.rf[28][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12398_ (.CLK(clknet_leaf_53_clk),
    .D(_00882_),
    .Q(\rvsingle.dp.rf.rf[28][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12399_ (.CLK(clknet_leaf_36_clk),
    .D(_00883_),
    .Q(\rvsingle.dp.rf.rf[28][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12400_ (.CLK(clknet_leaf_53_clk),
    .D(_00884_),
    .Q(\rvsingle.dp.rf.rf[28][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12401_ (.CLK(clknet_leaf_49_clk),
    .D(_00885_),
    .Q(\rvsingle.dp.rf.rf[28][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12402_ (.CLK(clknet_leaf_41_clk),
    .D(_00886_),
    .Q(\rvsingle.dp.rf.rf[28][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12403_ (.CLK(clknet_leaf_35_clk),
    .D(_00887_),
    .Q(\rvsingle.dp.rf.rf[28][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12404_ (.CLK(clknet_leaf_21_clk),
    .D(_00888_),
    .Q(\rvsingle.dp.rf.rf[28][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12405_ (.CLK(clknet_leaf_36_clk),
    .D(_00889_),
    .Q(\rvsingle.dp.rf.rf[28][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12406_ (.CLK(clknet_leaf_31_clk),
    .D(_00890_),
    .Q(\rvsingle.dp.rf.rf[28][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12407_ (.CLK(clknet_leaf_6_clk),
    .D(_00891_),
    .Q(\rvsingle.dp.rf.rf[28][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12408_ (.CLK(clknet_leaf_34_clk),
    .D(_00892_),
    .Q(\rvsingle.dp.rf.rf[28][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12409_ (.CLK(clknet_leaf_32_clk),
    .D(_00893_),
    .Q(\rvsingle.dp.rf.rf[28][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12410_ (.CLK(clknet_leaf_5_clk),
    .D(_00894_),
    .Q(\rvsingle.dp.rf.rf[28][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12411_ (.CLK(clknet_leaf_142_clk),
    .D(_00895_),
    .Q(\rvsingle.dp.rf.rf[28][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12412_ (.CLK(clknet_leaf_147_clk),
    .D(_00896_),
    .Q(\rvsingle.dp.rf.rf[28][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12413_ (.CLK(clknet_leaf_143_clk),
    .D(_00897_),
    .Q(\rvsingle.dp.rf.rf[28][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12414_ (.CLK(clknet_leaf_2_clk),
    .D(_00898_),
    .Q(\rvsingle.dp.rf.rf[28][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12415_ (.CLK(clknet_leaf_2_clk),
    .D(_00899_),
    .Q(\rvsingle.dp.rf.rf[28][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12416_ (.CLK(clknet_leaf_117_clk),
    .D(_00900_),
    .Q(\rvsingle.dp.rf.rf[28][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12417_ (.CLK(clknet_leaf_140_clk),
    .D(_00901_),
    .Q(\rvsingle.dp.rf.rf[28][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12418_ (.CLK(clknet_leaf_130_clk),
    .D(_00902_),
    .Q(\rvsingle.dp.rf.rf[28][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12419_ (.CLK(clknet_leaf_115_clk),
    .D(_00903_),
    .Q(\rvsingle.dp.rf.rf[28][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12420_ (.CLK(clknet_leaf_107_clk),
    .D(_00904_),
    .Q(\rvsingle.dp.rf.rf[28][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12421_ (.CLK(clknet_leaf_114_clk),
    .D(_00905_),
    .Q(\rvsingle.dp.rf.rf[28][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12422_ (.CLK(clknet_leaf_108_clk),
    .D(_00906_),
    .Q(\rvsingle.dp.rf.rf[28][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12423_ (.CLK(clknet_leaf_99_clk),
    .D(_00907_),
    .Q(\rvsingle.dp.rf.rf[28][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12424_ (.CLK(clknet_leaf_106_clk),
    .D(_00908_),
    .Q(\rvsingle.dp.rf.rf[28][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12425_ (.CLK(clknet_leaf_94_clk),
    .D(_00909_),
    .Q(\rvsingle.dp.rf.rf[28][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12426_ (.CLK(clknet_leaf_82_clk),
    .D(_00910_),
    .Q(\rvsingle.dp.rf.rf[28][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12427_ (.CLK(clknet_leaf_64_clk),
    .D(_00911_),
    .Q(\rvsingle.dp.rf.rf[27][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12428_ (.CLK(clknet_leaf_50_clk),
    .D(_00912_),
    .Q(\rvsingle.dp.rf.rf[27][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12429_ (.CLK(clknet_leaf_45_clk),
    .D(_00913_),
    .Q(\rvsingle.dp.rf.rf[27][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12430_ (.CLK(clknet_leaf_67_clk),
    .D(_00914_),
    .Q(\rvsingle.dp.rf.rf[27][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12431_ (.CLK(clknet_leaf_39_clk),
    .D(_00915_),
    .Q(\rvsingle.dp.rf.rf[27][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12432_ (.CLK(clknet_leaf_70_clk),
    .D(_00916_),
    .Q(\rvsingle.dp.rf.rf[27][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12433_ (.CLK(clknet_leaf_48_clk),
    .D(_00917_),
    .Q(\rvsingle.dp.rf.rf[27][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12434_ (.CLK(clknet_leaf_36_clk),
    .D(_00918_),
    .Q(\rvsingle.dp.rf.rf[27][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12435_ (.CLK(clknet_leaf_33_clk),
    .D(_00919_),
    .Q(\rvsingle.dp.rf.rf[27][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12436_ (.CLK(clknet_leaf_21_clk),
    .D(_00920_),
    .Q(\rvsingle.dp.rf.rf[27][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12437_ (.CLK(clknet_leaf_36_clk),
    .D(_00921_),
    .Q(\rvsingle.dp.rf.rf[27][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12438_ (.CLK(clknet_leaf_33_clk),
    .D(_00922_),
    .Q(\rvsingle.dp.rf.rf[27][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12439_ (.CLK(clknet_leaf_6_clk),
    .D(_00923_),
    .Q(\rvsingle.dp.rf.rf[27][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12440_ (.CLK(clknet_leaf_34_clk),
    .D(_00924_),
    .Q(\rvsingle.dp.rf.rf[27][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12441_ (.CLK(clknet_leaf_7_clk),
    .D(_00925_),
    .Q(\rvsingle.dp.rf.rf[27][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12442_ (.CLK(clknet_leaf_4_clk),
    .D(_00926_),
    .Q(\rvsingle.dp.rf.rf[27][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12443_ (.CLK(clknet_leaf_136_clk),
    .D(_00927_),
    .Q(\rvsingle.dp.rf.rf[27][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12444_ (.CLK(clknet_leaf_146_clk),
    .D(_00928_),
    .Q(\rvsingle.dp.rf.rf[27][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12445_ (.CLK(clknet_leaf_143_clk),
    .D(_00929_),
    .Q(\rvsingle.dp.rf.rf[27][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12446_ (.CLK(clknet_leaf_135_clk),
    .D(_00930_),
    .Q(\rvsingle.dp.rf.rf[27][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12447_ (.CLK(clknet_leaf_13_clk),
    .D(_00931_),
    .Q(\rvsingle.dp.rf.rf[27][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12448_ (.CLK(clknet_leaf_120_clk),
    .D(_00932_),
    .Q(\rvsingle.dp.rf.rf[27][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12449_ (.CLK(clknet_leaf_141_clk),
    .D(_00933_),
    .Q(\rvsingle.dp.rf.rf[27][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12450_ (.CLK(clknet_leaf_128_clk),
    .D(_00934_),
    .Q(\rvsingle.dp.rf.rf[27][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12451_ (.CLK(clknet_leaf_126_clk),
    .D(_00935_),
    .Q(\rvsingle.dp.rf.rf[27][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12452_ (.CLK(clknet_leaf_107_clk),
    .D(_00936_),
    .Q(\rvsingle.dp.rf.rf[27][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12453_ (.CLK(clknet_leaf_114_clk),
    .D(_00937_),
    .Q(\rvsingle.dp.rf.rf[27][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12454_ (.CLK(clknet_leaf_108_clk),
    .D(_00938_),
    .Q(\rvsingle.dp.rf.rf[27][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12455_ (.CLK(clknet_leaf_92_clk),
    .D(_00939_),
    .Q(\rvsingle.dp.rf.rf[27][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12456_ (.CLK(clknet_leaf_106_clk),
    .D(_00940_),
    .Q(\rvsingle.dp.rf.rf[27][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12457_ (.CLK(clknet_leaf_96_clk),
    .D(_00941_),
    .Q(\rvsingle.dp.rf.rf[27][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12458_ (.CLK(clknet_leaf_82_clk),
    .D(_00942_),
    .Q(\rvsingle.dp.rf.rf[27][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12459_ (.CLK(clknet_leaf_87_clk),
    .D(_00943_),
    .Q(\rvsingle.dp.rf.rf[26][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12460_ (.CLK(clknet_leaf_50_clk),
    .D(_00944_),
    .Q(\rvsingle.dp.rf.rf[26][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12461_ (.CLK(clknet_leaf_44_clk),
    .D(_00945_),
    .Q(\rvsingle.dp.rf.rf[26][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12462_ (.CLK(clknet_leaf_72_clk),
    .D(_00946_),
    .Q(\rvsingle.dp.rf.rf[26][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12463_ (.CLK(clknet_leaf_39_clk),
    .D(_00947_),
    .Q(\rvsingle.dp.rf.rf[26][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12464_ (.CLK(clknet_leaf_70_clk),
    .D(_00948_),
    .Q(\rvsingle.dp.rf.rf[26][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12465_ (.CLK(clknet_leaf_48_clk),
    .D(_00949_),
    .Q(\rvsingle.dp.rf.rf[26][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12466_ (.CLK(clknet_leaf_27_clk),
    .D(_00950_),
    .Q(\rvsingle.dp.rf.rf[26][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12467_ (.CLK(clknet_leaf_29_clk),
    .D(_00951_),
    .Q(\rvsingle.dp.rf.rf[26][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12468_ (.CLK(clknet_leaf_20_clk),
    .D(_00952_),
    .Q(\rvsingle.dp.rf.rf[26][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12469_ (.CLK(clknet_leaf_27_clk),
    .D(_00953_),
    .Q(\rvsingle.dp.rf.rf[26][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12470_ (.CLK(clknet_leaf_31_clk),
    .D(_00954_),
    .Q(\rvsingle.dp.rf.rf[26][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12471_ (.CLK(clknet_leaf_6_clk),
    .D(_00955_),
    .Q(\rvsingle.dp.rf.rf[26][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12472_ (.CLK(clknet_leaf_34_clk),
    .D(_00956_),
    .Q(\rvsingle.dp.rf.rf[26][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12473_ (.CLK(clknet_leaf_8_clk),
    .D(_00957_),
    .Q(\rvsingle.dp.rf.rf[26][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12474_ (.CLK(clknet_leaf_5_clk),
    .D(_00958_),
    .Q(\rvsingle.dp.rf.rf[26][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12475_ (.CLK(clknet_leaf_136_clk),
    .D(_00959_),
    .Q(\rvsingle.dp.rf.rf[26][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12476_ (.CLK(clknet_leaf_151_clk),
    .D(_00960_),
    .Q(\rvsingle.dp.rf.rf[26][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12477_ (.CLK(clknet_leaf_146_clk),
    .D(_00961_),
    .Q(\rvsingle.dp.rf.rf[26][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12478_ (.CLK(clknet_leaf_150_clk),
    .D(_00962_),
    .Q(\rvsingle.dp.rf.rf[26][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12479_ (.CLK(clknet_leaf_1_clk),
    .D(_00963_),
    .Q(\rvsingle.dp.rf.rf[26][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12480_ (.CLK(clknet_leaf_118_clk),
    .D(_00964_),
    .Q(\rvsingle.dp.rf.rf[26][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12481_ (.CLK(clknet_leaf_140_clk),
    .D(_00965_),
    .Q(\rvsingle.dp.rf.rf[26][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12482_ (.CLK(clknet_leaf_128_clk),
    .D(_00966_),
    .Q(\rvsingle.dp.rf.rf[26][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12483_ (.CLK(clknet_leaf_126_clk),
    .D(_00967_),
    .Q(\rvsingle.dp.rf.rf[26][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12484_ (.CLK(clknet_leaf_109_clk),
    .D(_00968_),
    .Q(\rvsingle.dp.rf.rf[26][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12485_ (.CLK(clknet_leaf_114_clk),
    .D(_00969_),
    .Q(\rvsingle.dp.rf.rf[26][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12486_ (.CLK(clknet_leaf_108_clk),
    .D(_00970_),
    .Q(\rvsingle.dp.rf.rf[26][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12487_ (.CLK(clknet_leaf_101_clk),
    .D(_00971_),
    .Q(\rvsingle.dp.rf.rf[26][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12488_ (.CLK(clknet_leaf_106_clk),
    .D(_00972_),
    .Q(\rvsingle.dp.rf.rf[26][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12489_ (.CLK(clknet_leaf_96_clk),
    .D(_00973_),
    .Q(\rvsingle.dp.rf.rf[26][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12490_ (.CLK(clknet_leaf_82_clk),
    .D(_00974_),
    .Q(\rvsingle.dp.rf.rf[26][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12491_ (.CLK(clknet_leaf_64_clk),
    .D(_00975_),
    .Q(\rvsingle.dp.rf.rf[25][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12492_ (.CLK(clknet_leaf_50_clk),
    .D(_00976_),
    .Q(\rvsingle.dp.rf.rf[25][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12493_ (.CLK(clknet_leaf_44_clk),
    .D(_00977_),
    .Q(\rvsingle.dp.rf.rf[25][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12494_ (.CLK(clknet_leaf_67_clk),
    .D(_00978_),
    .Q(\rvsingle.dp.rf.rf[25][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12495_ (.CLK(clknet_leaf_39_clk),
    .D(_00979_),
    .Q(\rvsingle.dp.rf.rf[25][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12496_ (.CLK(clknet_leaf_70_clk),
    .D(_00980_),
    .Q(\rvsingle.dp.rf.rf[25][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12497_ (.CLK(clknet_leaf_48_clk),
    .D(_00981_),
    .Q(\rvsingle.dp.rf.rf[25][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12498_ (.CLK(clknet_leaf_36_clk),
    .D(_00982_),
    .Q(\rvsingle.dp.rf.rf[25][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12499_ (.CLK(clknet_leaf_33_clk),
    .D(_00983_),
    .Q(\rvsingle.dp.rf.rf[25][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12500_ (.CLK(clknet_leaf_21_clk),
    .D(_00984_),
    .Q(\rvsingle.dp.rf.rf[25][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12501_ (.CLK(clknet_leaf_36_clk),
    .D(_00985_),
    .Q(\rvsingle.dp.rf.rf[25][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12502_ (.CLK(clknet_leaf_34_clk),
    .D(_00986_),
    .Q(\rvsingle.dp.rf.rf[25][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12503_ (.CLK(clknet_leaf_6_clk),
    .D(_00987_),
    .Q(\rvsingle.dp.rf.rf[25][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12504_ (.CLK(clknet_leaf_34_clk),
    .D(_00988_),
    .Q(\rvsingle.dp.rf.rf[25][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12505_ (.CLK(clknet_leaf_7_clk),
    .D(_00989_),
    .Q(\rvsingle.dp.rf.rf[25][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12506_ (.CLK(clknet_leaf_4_clk),
    .D(_00990_),
    .Q(\rvsingle.dp.rf.rf[25][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12507_ (.CLK(clknet_leaf_136_clk),
    .D(_00991_),
    .Q(\rvsingle.dp.rf.rf[25][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12508_ (.CLK(clknet_leaf_146_clk),
    .D(_00992_),
    .Q(\rvsingle.dp.rf.rf[25][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12509_ (.CLK(clknet_leaf_143_clk),
    .D(_00993_),
    .Q(\rvsingle.dp.rf.rf[25][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12510_ (.CLK(clknet_leaf_135_clk),
    .D(_00994_),
    .Q(\rvsingle.dp.rf.rf[25][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12511_ (.CLK(clknet_leaf_13_clk),
    .D(_00995_),
    .Q(\rvsingle.dp.rf.rf[25][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12512_ (.CLK(clknet_leaf_119_clk),
    .D(_00996_),
    .Q(\rvsingle.dp.rf.rf[25][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12513_ (.CLK(clknet_leaf_139_clk),
    .D(_00997_),
    .Q(\rvsingle.dp.rf.rf[25][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12514_ (.CLK(clknet_leaf_128_clk),
    .D(_00998_),
    .Q(\rvsingle.dp.rf.rf[25][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12515_ (.CLK(clknet_leaf_127_clk),
    .D(_00999_),
    .Q(\rvsingle.dp.rf.rf[25][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12516_ (.CLK(clknet_leaf_108_clk),
    .D(_01000_),
    .Q(\rvsingle.dp.rf.rf[25][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12517_ (.CLK(clknet_leaf_115_clk),
    .D(_01001_),
    .Q(\rvsingle.dp.rf.rf[25][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12518_ (.CLK(clknet_leaf_108_clk),
    .D(_01002_),
    .Q(\rvsingle.dp.rf.rf[25][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12519_ (.CLK(clknet_leaf_100_clk),
    .D(_01003_),
    .Q(\rvsingle.dp.rf.rf[25][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12520_ (.CLK(clknet_leaf_106_clk),
    .D(_01004_),
    .Q(\rvsingle.dp.rf.rf[25][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12521_ (.CLK(clknet_leaf_96_clk),
    .D(_01005_),
    .Q(\rvsingle.dp.rf.rf[25][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12522_ (.CLK(clknet_leaf_83_clk),
    .D(_01006_),
    .Q(\rvsingle.dp.rf.rf[25][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12523_ (.CLK(clknet_leaf_86_clk),
    .D(_01007_),
    .Q(\rvsingle.dp.rf.rf[24][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12524_ (.CLK(clknet_leaf_50_clk),
    .D(_01008_),
    .Q(\rvsingle.dp.rf.rf[24][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12525_ (.CLK(clknet_leaf_44_clk),
    .D(_01009_),
    .Q(\rvsingle.dp.rf.rf[24][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12526_ (.CLK(clknet_leaf_72_clk),
    .D(_01010_),
    .Q(\rvsingle.dp.rf.rf[24][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12527_ (.CLK(clknet_leaf_39_clk),
    .D(_01011_),
    .Q(\rvsingle.dp.rf.rf[24][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12528_ (.CLK(clknet_leaf_70_clk),
    .D(_01012_),
    .Q(\rvsingle.dp.rf.rf[24][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12529_ (.CLK(clknet_leaf_49_clk),
    .D(_01013_),
    .Q(\rvsingle.dp.rf.rf[24][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12530_ (.CLK(clknet_leaf_35_clk),
    .D(_01014_),
    .Q(\rvsingle.dp.rf.rf[24][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12531_ (.CLK(clknet_leaf_32_clk),
    .D(_01015_),
    .Q(\rvsingle.dp.rf.rf[24][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12532_ (.CLK(clknet_leaf_62_clk),
    .D(_01016_),
    .Q(\rvsingle.dp.rf.rf[24][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12533_ (.CLK(clknet_leaf_36_clk),
    .D(_01017_),
    .Q(\rvsingle.dp.rf.rf[24][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12534_ (.CLK(clknet_leaf_35_clk),
    .D(_01018_),
    .Q(\rvsingle.dp.rf.rf[24][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12535_ (.CLK(clknet_leaf_15_clk),
    .D(_01019_),
    .Q(\rvsingle.dp.rf.rf[24][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12536_ (.CLK(clknet_leaf_34_clk),
    .D(_01020_),
    .Q(\rvsingle.dp.rf.rf[24][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12537_ (.CLK(clknet_leaf_7_clk),
    .D(_01021_),
    .Q(\rvsingle.dp.rf.rf[24][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12538_ (.CLK(clknet_leaf_4_clk),
    .D(_01022_),
    .Q(\rvsingle.dp.rf.rf[24][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12539_ (.CLK(clknet_leaf_145_clk),
    .D(_01023_),
    .Q(\rvsingle.dp.rf.rf[24][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12540_ (.CLK(clknet_leaf_151_clk),
    .D(_01024_),
    .Q(\rvsingle.dp.rf.rf[24][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12541_ (.CLK(clknet_leaf_143_clk),
    .D(_01025_),
    .Q(\rvsingle.dp.rf.rf[24][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12542_ (.CLK(clknet_leaf_0_clk),
    .D(_01026_),
    .Q(\rvsingle.dp.rf.rf[24][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12543_ (.CLK(clknet_leaf_1_clk),
    .D(_01027_),
    .Q(\rvsingle.dp.rf.rf[24][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12544_ (.CLK(clknet_leaf_117_clk),
    .D(_01028_),
    .Q(\rvsingle.dp.rf.rf[24][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12545_ (.CLK(clknet_leaf_141_clk),
    .D(_01029_),
    .Q(\rvsingle.dp.rf.rf[24][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12546_ (.CLK(clknet_leaf_126_clk),
    .D(_01030_),
    .Q(\rvsingle.dp.rf.rf[24][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12547_ (.CLK(clknet_leaf_127_clk),
    .D(_01031_),
    .Q(\rvsingle.dp.rf.rf[24][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12548_ (.CLK(clknet_leaf_107_clk),
    .D(_01032_),
    .Q(\rvsingle.dp.rf.rf[24][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12549_ (.CLK(clknet_leaf_114_clk),
    .D(_01033_),
    .Q(\rvsingle.dp.rf.rf[24][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12550_ (.CLK(clknet_leaf_108_clk),
    .D(_01034_),
    .Q(\rvsingle.dp.rf.rf[24][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12551_ (.CLK(clknet_leaf_127_clk),
    .D(_01035_),
    .Q(\rvsingle.dp.rf.rf[24][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12552_ (.CLK(clknet_leaf_106_clk),
    .D(_01036_),
    .Q(\rvsingle.dp.rf.rf[24][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12553_ (.CLK(clknet_leaf_96_clk),
    .D(_01037_),
    .Q(\rvsingle.dp.rf.rf[24][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12554_ (.CLK(clknet_leaf_84_clk),
    .D(_01038_),
    .Q(\rvsingle.dp.rf.rf[24][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12555_ (.CLK(clknet_leaf_88_clk),
    .D(_01039_),
    .Q(\rvsingle.dp.rf.rf[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12556_ (.CLK(clknet_leaf_51_clk),
    .D(_01040_),
    .Q(\rvsingle.dp.rf.rf[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12557_ (.CLK(clknet_leaf_43_clk),
    .D(_01041_),
    .Q(\rvsingle.dp.rf.rf[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12558_ (.CLK(clknet_leaf_68_clk),
    .D(_01042_),
    .Q(\rvsingle.dp.rf.rf[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12559_ (.CLK(clknet_leaf_57_clk),
    .D(_01043_),
    .Q(\rvsingle.dp.rf.rf[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12560_ (.CLK(clknet_leaf_68_clk),
    .D(_01044_),
    .Q(\rvsingle.dp.rf.rf[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12561_ (.CLK(clknet_leaf_48_clk),
    .D(_01045_),
    .Q(\rvsingle.dp.rf.rf[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12562_ (.CLK(clknet_leaf_59_clk),
    .D(_01046_),
    .Q(\rvsingle.dp.rf.rf[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12563_ (.CLK(clknet_4_8_0_clk),
    .D(_01047_),
    .Q(\rvsingle.dp.rf.rf[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12564_ (.CLK(clknet_leaf_21_clk),
    .D(_01048_),
    .Q(\rvsingle.dp.rf.rf[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12565_ (.CLK(clknet_leaf_64_clk),
    .D(_01049_),
    .Q(\rvsingle.dp.rf.rf[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12566_ (.CLK(clknet_leaf_25_clk),
    .D(_01050_),
    .Q(\rvsingle.dp.rf.rf[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12567_ (.CLK(clknet_leaf_16_clk),
    .D(_01051_),
    .Q(\rvsingle.dp.rf.rf[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12568_ (.CLK(clknet_leaf_22_clk),
    .D(_01052_),
    .Q(\rvsingle.dp.rf.rf[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12569_ (.CLK(clknet_leaf_16_clk),
    .D(_01053_),
    .Q(\rvsingle.dp.rf.rf[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12570_ (.CLK(clknet_leaf_5_clk),
    .D(_01054_),
    .Q(\rvsingle.dp.rf.rf[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12571_ (.CLK(clknet_leaf_136_clk),
    .D(_01055_),
    .Q(\rvsingle.dp.rf.rf[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12572_ (.CLK(clknet_leaf_150_clk),
    .D(_01056_),
    .Q(\rvsingle.dp.rf.rf[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12573_ (.CLK(clknet_leaf_133_clk),
    .D(_01057_),
    .Q(\rvsingle.dp.rf.rf[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12574_ (.CLK(clknet_leaf_146_clk),
    .D(_00032_),
    .Q(\rvsingle.dp.rf.rf[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12575_ (.CLK(clknet_leaf_2_clk),
    .D(_00033_),
    .Q(\rvsingle.dp.rf.rf[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12576_ (.CLK(clknet_leaf_120_clk),
    .D(_00034_),
    .Q(\rvsingle.dp.rf.rf[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12577_ (.CLK(clknet_leaf_130_clk),
    .D(_00035_),
    .Q(\rvsingle.dp.rf.rf[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12578_ (.CLK(clknet_leaf_128_clk),
    .D(_00036_),
    .Q(\rvsingle.dp.rf.rf[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12579_ (.CLK(clknet_leaf_121_clk),
    .D(_00037_),
    .Q(\rvsingle.dp.rf.rf[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12580_ (.CLK(clknet_leaf_123_clk),
    .D(_00038_),
    .Q(\rvsingle.dp.rf.rf[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12581_ (.CLK(clknet_leaf_123_clk),
    .D(_00039_),
    .Q(\rvsingle.dp.rf.rf[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12582_ (.CLK(clknet_leaf_122_clk),
    .D(_00040_),
    .Q(\rvsingle.dp.rf.rf[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12583_ (.CLK(clknet_leaf_101_clk),
    .D(_00041_),
    .Q(\rvsingle.dp.rf.rf[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12584_ (.CLK(clknet_leaf_123_clk),
    .D(_00042_),
    .Q(\rvsingle.dp.rf.rf[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12585_ (.CLK(clknet_leaf_97_clk),
    .D(_00043_),
    .Q(\rvsingle.dp.rf.rf[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12586_ (.CLK(clknet_leaf_83_clk),
    .D(_00044_),
    .Q(\rvsingle.dp.rf.rf[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12587_ (.CLK(clknet_leaf_87_clk),
    .D(_00045_),
    .Q(\rvsingle.dp.rf.rf[22][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12588_ (.CLK(clknet_leaf_49_clk),
    .D(_00046_),
    .Q(\rvsingle.dp.rf.rf[22][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12589_ (.CLK(clknet_leaf_44_clk),
    .D(_00047_),
    .Q(\rvsingle.dp.rf.rf[22][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12590_ (.CLK(clknet_leaf_71_clk),
    .D(_00048_),
    .Q(\rvsingle.dp.rf.rf[22][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12591_ (.CLK(clknet_leaf_37_clk),
    .D(_00049_),
    .Q(\rvsingle.dp.rf.rf[22][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12592_ (.CLK(clknet_leaf_71_clk),
    .D(_00050_),
    .Q(\rvsingle.dp.rf.rf[22][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12593_ (.CLK(clknet_leaf_49_clk),
    .D(_00051_),
    .Q(\rvsingle.dp.rf.rf[22][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12594_ (.CLK(clknet_leaf_39_clk),
    .D(_00052_),
    .Q(\rvsingle.dp.rf.rf[22][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12595_ (.CLK(clknet_leaf_35_clk),
    .D(_00053_),
    .Q(\rvsingle.dp.rf.rf[22][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12596_ (.CLK(clknet_leaf_58_clk),
    .D(_00054_),
    .Q(\rvsingle.dp.rf.rf[22][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12597_ (.CLK(clknet_leaf_37_clk),
    .D(_00055_),
    .Q(\rvsingle.dp.rf.rf[22][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12598_ (.CLK(clknet_leaf_33_clk),
    .D(_00056_),
    .Q(\rvsingle.dp.rf.rf[22][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12599_ (.CLK(clknet_leaf_7_clk),
    .D(_00057_),
    .Q(\rvsingle.dp.rf.rf[22][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12600_ (.CLK(clknet_leaf_33_clk),
    .D(_00058_),
    .Q(\rvsingle.dp.rf.rf[22][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12601_ (.CLK(clknet_leaf_7_clk),
    .D(_00059_),
    .Q(\rvsingle.dp.rf.rf[22][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12602_ (.CLK(clknet_leaf_3_clk),
    .D(_00060_),
    .Q(\rvsingle.dp.rf.rf[22][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12603_ (.CLK(clknet_leaf_142_clk),
    .D(_00061_),
    .Q(\rvsingle.dp.rf.rf[22][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12604_ (.CLK(clknet_leaf_149_clk),
    .D(_00062_),
    .Q(\rvsingle.dp.rf.rf[22][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12605_ (.CLK(clknet_leaf_143_clk),
    .D(_00063_),
    .Q(\rvsingle.dp.rf.rf[22][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12606_ (.CLK(clknet_leaf_150_clk),
    .D(_00064_),
    .Q(\rvsingle.dp.rf.rf[22][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12607_ (.CLK(clknet_leaf_0_clk),
    .D(_00065_),
    .Q(\rvsingle.dp.rf.rf[22][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12608_ (.CLK(clknet_leaf_118_clk),
    .D(_00066_),
    .Q(\rvsingle.dp.rf.rf[22][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12609_ (.CLK(clknet_leaf_140_clk),
    .D(_00067_),
    .Q(\rvsingle.dp.rf.rf[22][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12610_ (.CLK(clknet_leaf_128_clk),
    .D(_00068_),
    .Q(\rvsingle.dp.rf.rf[22][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12611_ (.CLK(clknet_leaf_115_clk),
    .D(_00069_),
    .Q(\rvsingle.dp.rf.rf[22][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12612_ (.CLK(clknet_leaf_107_clk),
    .D(_00070_),
    .Q(\rvsingle.dp.rf.rf[22][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12613_ (.CLK(clknet_leaf_115_clk),
    .D(_00071_),
    .Q(\rvsingle.dp.rf.rf[22][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12614_ (.CLK(clknet_leaf_113_clk),
    .D(_00072_),
    .Q(\rvsingle.dp.rf.rf[22][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12615_ (.CLK(clknet_leaf_104_clk),
    .D(_00073_),
    .Q(\rvsingle.dp.rf.rf[22][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12616_ (.CLK(clknet_leaf_106_clk),
    .D(_00074_),
    .Q(\rvsingle.dp.rf.rf[22][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12617_ (.CLK(clknet_leaf_95_clk),
    .D(_00075_),
    .Q(\rvsingle.dp.rf.rf[22][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12618_ (.CLK(clknet_leaf_83_clk),
    .D(_00076_),
    .Q(\rvsingle.dp.rf.rf[22][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12619_ (.CLK(clknet_leaf_64_clk),
    .D(_00077_),
    .Q(\rvsingle.dp.rf.rf[21][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12620_ (.CLK(clknet_leaf_50_clk),
    .D(_00078_),
    .Q(\rvsingle.dp.rf.rf[21][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12621_ (.CLK(clknet_leaf_43_clk),
    .D(_00079_),
    .Q(\rvsingle.dp.rf.rf[21][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12622_ (.CLK(clknet_leaf_71_clk),
    .D(_00080_),
    .Q(\rvsingle.dp.rf.rf[21][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12623_ (.CLK(clknet_leaf_36_clk),
    .D(_00081_),
    .Q(\rvsingle.dp.rf.rf[21][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12624_ (.CLK(clknet_leaf_70_clk),
    .D(_00082_),
    .Q(\rvsingle.dp.rf.rf[21][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12625_ (.CLK(clknet_leaf_48_clk),
    .D(_00083_),
    .Q(\rvsingle.dp.rf.rf[21][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12626_ (.CLK(clknet_leaf_41_clk),
    .D(_00084_),
    .Q(\rvsingle.dp.rf.rf[21][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12627_ (.CLK(clknet_leaf_35_clk),
    .D(_00085_),
    .Q(\rvsingle.dp.rf.rf[21][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12628_ (.CLK(clknet_leaf_59_clk),
    .D(_00086_),
    .Q(\rvsingle.dp.rf.rf[21][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12629_ (.CLK(clknet_leaf_36_clk),
    .D(_00087_),
    .Q(\rvsingle.dp.rf.rf[21][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12630_ (.CLK(clknet_leaf_33_clk),
    .D(_00088_),
    .Q(\rvsingle.dp.rf.rf[21][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12631_ (.CLK(clknet_leaf_6_clk),
    .D(_00089_),
    .Q(\rvsingle.dp.rf.rf[21][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12632_ (.CLK(clknet_leaf_33_clk),
    .D(_00090_),
    .Q(\rvsingle.dp.rf.rf[21][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12633_ (.CLK(clknet_leaf_8_clk),
    .D(_00091_),
    .Q(\rvsingle.dp.rf.rf[21][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12634_ (.CLK(clknet_leaf_3_clk),
    .D(_00092_),
    .Q(\rvsingle.dp.rf.rf[21][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12635_ (.CLK(clknet_leaf_142_clk),
    .D(_00093_),
    .Q(\rvsingle.dp.rf.rf[21][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12636_ (.CLK(clknet_leaf_151_clk),
    .D(_00094_),
    .Q(\rvsingle.dp.rf.rf[21][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12637_ (.CLK(clknet_leaf_144_clk),
    .D(_00095_),
    .Q(\rvsingle.dp.rf.rf[21][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12638_ (.CLK(clknet_leaf_150_clk),
    .D(_00096_),
    .Q(\rvsingle.dp.rf.rf[21][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12639_ (.CLK(clknet_leaf_2_clk),
    .D(_00097_),
    .Q(\rvsingle.dp.rf.rf[21][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12640_ (.CLK(clknet_leaf_118_clk),
    .D(_00098_),
    .Q(\rvsingle.dp.rf.rf[21][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12641_ (.CLK(clknet_leaf_140_clk),
    .D(_00099_),
    .Q(\rvsingle.dp.rf.rf[21][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12642_ (.CLK(clknet_leaf_128_clk),
    .D(_00100_),
    .Q(\rvsingle.dp.rf.rf[21][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12643_ (.CLK(clknet_leaf_115_clk),
    .D(_00101_),
    .Q(\rvsingle.dp.rf.rf[21][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12644_ (.CLK(clknet_leaf_107_clk),
    .D(_00102_),
    .Q(\rvsingle.dp.rf.rf[21][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12645_ (.CLK(clknet_leaf_115_clk),
    .D(_00103_),
    .Q(\rvsingle.dp.rf.rf[21][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12646_ (.CLK(clknet_leaf_113_clk),
    .D(_00104_),
    .Q(\rvsingle.dp.rf.rf[21][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12647_ (.CLK(clknet_leaf_104_clk),
    .D(_00105_),
    .Q(\rvsingle.dp.rf.rf[21][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12648_ (.CLK(clknet_leaf_105_clk),
    .D(_00106_),
    .Q(\rvsingle.dp.rf.rf[21][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12649_ (.CLK(clknet_leaf_95_clk),
    .D(_00107_),
    .Q(\rvsingle.dp.rf.rf[21][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12650_ (.CLK(clknet_leaf_82_clk),
    .D(_00108_),
    .Q(\rvsingle.dp.rf.rf[21][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12651_ (.CLK(clknet_leaf_64_clk),
    .D(_00109_),
    .Q(\rvsingle.dp.rf.rf[20][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12652_ (.CLK(clknet_leaf_49_clk),
    .D(_00110_),
    .Q(\rvsingle.dp.rf.rf[20][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12653_ (.CLK(clknet_leaf_43_clk),
    .D(_00111_),
    .Q(\rvsingle.dp.rf.rf[20][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12654_ (.CLK(clknet_leaf_72_clk),
    .D(_00112_),
    .Q(\rvsingle.dp.rf.rf[20][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12655_ (.CLK(clknet_leaf_36_clk),
    .D(_00113_),
    .Q(\rvsingle.dp.rf.rf[20][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12656_ (.CLK(clknet_leaf_72_clk),
    .D(_00114_),
    .Q(\rvsingle.dp.rf.rf[20][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12657_ (.CLK(clknet_leaf_49_clk),
    .D(_00115_),
    .Q(\rvsingle.dp.rf.rf[20][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12658_ (.CLK(clknet_leaf_41_clk),
    .D(_00116_),
    .Q(\rvsingle.dp.rf.rf[20][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12659_ (.CLK(clknet_leaf_35_clk),
    .D(_00117_),
    .Q(\rvsingle.dp.rf.rf[20][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12660_ (.CLK(clknet_leaf_59_clk),
    .D(_00118_),
    .Q(\rvsingle.dp.rf.rf[20][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12661_ (.CLK(clknet_leaf_36_clk),
    .D(_00119_),
    .Q(\rvsingle.dp.rf.rf[20][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12662_ (.CLK(clknet_leaf_33_clk),
    .D(_00120_),
    .Q(\rvsingle.dp.rf.rf[20][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12663_ (.CLK(clknet_leaf_7_clk),
    .D(_00121_),
    .Q(\rvsingle.dp.rf.rf[20][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12664_ (.CLK(clknet_leaf_33_clk),
    .D(_00122_),
    .Q(\rvsingle.dp.rf.rf[20][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12665_ (.CLK(clknet_leaf_8_clk),
    .D(_00123_),
    .Q(\rvsingle.dp.rf.rf[20][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12666_ (.CLK(clknet_leaf_3_clk),
    .D(_00124_),
    .Q(\rvsingle.dp.rf.rf[20][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12667_ (.CLK(clknet_leaf_141_clk),
    .D(_00125_),
    .Q(\rvsingle.dp.rf.rf[20][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12668_ (.CLK(clknet_leaf_151_clk),
    .D(_00126_),
    .Q(\rvsingle.dp.rf.rf[20][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12669_ (.CLK(clknet_leaf_143_clk),
    .D(_00127_),
    .Q(\rvsingle.dp.rf.rf[20][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12670_ (.CLK(clknet_leaf_150_clk),
    .D(_00128_),
    .Q(\rvsingle.dp.rf.rf[20][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12671_ (.CLK(clknet_leaf_2_clk),
    .D(_00129_),
    .Q(\rvsingle.dp.rf.rf[20][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12672_ (.CLK(clknet_leaf_117_clk),
    .D(_00130_),
    .Q(\rvsingle.dp.rf.rf[20][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12673_ (.CLK(clknet_leaf_140_clk),
    .D(_00131_),
    .Q(\rvsingle.dp.rf.rf[20][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12674_ (.CLK(clknet_leaf_128_clk),
    .D(_00132_),
    .Q(\rvsingle.dp.rf.rf[20][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12675_ (.CLK(clknet_leaf_115_clk),
    .D(_00133_),
    .Q(\rvsingle.dp.rf.rf[20][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12676_ (.CLK(clknet_leaf_107_clk),
    .D(_00134_),
    .Q(\rvsingle.dp.rf.rf[20][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12677_ (.CLK(clknet_leaf_114_clk),
    .D(_00135_),
    .Q(\rvsingle.dp.rf.rf[20][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12678_ (.CLK(clknet_leaf_113_clk),
    .D(_00136_),
    .Q(\rvsingle.dp.rf.rf[20][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12679_ (.CLK(clknet_leaf_104_clk),
    .D(_00137_),
    .Q(\rvsingle.dp.rf.rf[20][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12680_ (.CLK(clknet_leaf_105_clk),
    .D(_00138_),
    .Q(\rvsingle.dp.rf.rf[20][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12681_ (.CLK(clknet_leaf_95_clk),
    .D(_00139_),
    .Q(\rvsingle.dp.rf.rf[20][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12682_ (.CLK(clknet_leaf_82_clk),
    .D(_00140_),
    .Q(\rvsingle.dp.rf.rf[20][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12683_ (.CLK(clknet_leaf_88_clk),
    .D(_00141_),
    .Q(\rvsingle.dp.rf.rf[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12684_ (.CLK(clknet_leaf_54_clk),
    .D(_00142_),
    .Q(\rvsingle.dp.rf.rf[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12685_ (.CLK(clknet_leaf_45_clk),
    .D(_00143_),
    .Q(\rvsingle.dp.rf.rf[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12686_ (.CLK(clknet_leaf_67_clk),
    .D(_00144_),
    .Q(\rvsingle.dp.rf.rf[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12687_ (.CLK(clknet_leaf_59_clk),
    .D(_00145_),
    .Q(\rvsingle.dp.rf.rf[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12688_ (.CLK(clknet_leaf_67_clk),
    .D(_00146_),
    .Q(\rvsingle.dp.rf.rf[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12689_ (.CLK(clknet_leaf_67_clk),
    .D(_00147_),
    .Q(\rvsingle.dp.rf.rf[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12690_ (.CLK(clknet_leaf_27_clk),
    .D(_00148_),
    .Q(\rvsingle.dp.rf.rf[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12691_ (.CLK(clknet_leaf_28_clk),
    .D(_00149_),
    .Q(\rvsingle.dp.rf.rf[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12692_ (.CLK(clknet_leaf_62_clk),
    .D(_00150_),
    .Q(\rvsingle.dp.rf.rf[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12693_ (.CLK(clknet_leaf_60_clk),
    .D(_00151_),
    .Q(\rvsingle.dp.rf.rf[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12694_ (.CLK(clknet_leaf_26_clk),
    .D(_00152_),
    .Q(\rvsingle.dp.rf.rf[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12695_ (.CLK(clknet_leaf_18_clk),
    .D(_00153_),
    .Q(\rvsingle.dp.rf.rf[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12696_ (.CLK(clknet_leaf_19_clk),
    .D(_00154_),
    .Q(\rvsingle.dp.rf.rf[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12697_ (.CLK(clknet_leaf_23_clk),
    .D(_00155_),
    .Q(\rvsingle.dp.rf.rf[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12698_ (.CLK(clknet_leaf_15_clk),
    .D(_00156_),
    .Q(\rvsingle.dp.rf.rf[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12699_ (.CLK(clknet_leaf_137_clk),
    .D(_00157_),
    .Q(\rvsingle.dp.rf.rf[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12700_ (.CLK(clknet_leaf_146_clk),
    .D(_00158_),
    .Q(\rvsingle.dp.rf.rf[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12701_ (.CLK(clknet_leaf_136_clk),
    .D(_00159_),
    .Q(\rvsingle.dp.rf.rf[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12702_ (.CLK(clknet_leaf_133_clk),
    .D(_00160_),
    .Q(\rvsingle.dp.rf.rf[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12703_ (.CLK(clknet_leaf_131_clk),
    .D(_00161_),
    .Q(\rvsingle.dp.rf.rf[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12704_ (.CLK(clknet_leaf_120_clk),
    .D(_00162_),
    .Q(\rvsingle.dp.rf.rf[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12705_ (.CLK(clknet_leaf_125_clk),
    .D(_00163_),
    .Q(\rvsingle.dp.rf.rf[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12706_ (.CLK(clknet_leaf_131_clk),
    .D(_00164_),
    .Q(\rvsingle.dp.rf.rf[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12707_ (.CLK(clknet_leaf_124_clk),
    .D(_00165_),
    .Q(\rvsingle.dp.rf.rf[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12708_ (.CLK(clknet_leaf_124_clk),
    .D(_00166_),
    .Q(\rvsingle.dp.rf.rf[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12709_ (.CLK(clknet_leaf_110_clk),
    .D(_00167_),
    .Q(\rvsingle.dp.rf.rf[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12710_ (.CLK(clknet_leaf_115_clk),
    .D(_00168_),
    .Q(\rvsingle.dp.rf.rf[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12711_ (.CLK(clknet_leaf_98_clk),
    .D(_00169_),
    .Q(\rvsingle.dp.rf.rf[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12712_ (.CLK(clknet_leaf_104_clk),
    .D(_00170_),
    .Q(\rvsingle.dp.rf.rf[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12713_ (.CLK(clknet_leaf_127_clk),
    .D(_00171_),
    .Q(\rvsingle.dp.rf.rf[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12714_ (.CLK(clknet_leaf_95_clk),
    .D(_00172_),
    .Q(\rvsingle.dp.rf.rf[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12715_ (.CLK(clknet_leaf_86_clk),
    .D(_00173_),
    .Q(\rvsingle.dp.rf.rf[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12716_ (.CLK(clknet_leaf_50_clk),
    .D(_00174_),
    .Q(\rvsingle.dp.rf.rf[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12717_ (.CLK(clknet_leaf_45_clk),
    .D(_00175_),
    .Q(\rvsingle.dp.rf.rf[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12718_ (.CLK(clknet_leaf_71_clk),
    .D(_00176_),
    .Q(\rvsingle.dp.rf.rf[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12719_ (.CLK(clknet_leaf_27_clk),
    .D(_00177_),
    .Q(\rvsingle.dp.rf.rf[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12720_ (.CLK(clknet_leaf_52_clk),
    .D(_00178_),
    .Q(\rvsingle.dp.rf.rf[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12721_ (.CLK(clknet_leaf_49_clk),
    .D(_00179_),
    .Q(\rvsingle.dp.rf.rf[18][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12722_ (.CLK(clknet_leaf_47_clk),
    .D(_00180_),
    .Q(\rvsingle.dp.rf.rf[18][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12723_ (.CLK(clknet_leaf_27_clk),
    .D(_00181_),
    .Q(\rvsingle.dp.rf.rf[18][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12724_ (.CLK(clknet_leaf_61_clk),
    .D(_00182_),
    .Q(\rvsingle.dp.rf.rf[18][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12725_ (.CLK(clknet_leaf_58_clk),
    .D(_00183_),
    .Q(\rvsingle.dp.rf.rf[18][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12726_ (.CLK(clknet_leaf_32_clk),
    .D(_00184_),
    .Q(\rvsingle.dp.rf.rf[18][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12727_ (.CLK(clknet_leaf_6_clk),
    .D(_00185_),
    .Q(\rvsingle.dp.rf.rf[18][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12728_ (.CLK(clknet_leaf_32_clk),
    .D(_00186_),
    .Q(\rvsingle.dp.rf.rf[18][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12729_ (.CLK(clknet_leaf_8_clk),
    .D(_00187_),
    .Q(\rvsingle.dp.rf.rf[18][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12730_ (.CLK(clknet_leaf_4_clk),
    .D(_00188_),
    .Q(\rvsingle.dp.rf.rf[18][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12731_ (.CLK(clknet_leaf_141_clk),
    .D(_00189_),
    .Q(\rvsingle.dp.rf.rf[18][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12732_ (.CLK(clknet_leaf_147_clk),
    .D(_00190_),
    .Q(\rvsingle.dp.rf.rf[18][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12733_ (.CLK(clknet_leaf_143_clk),
    .D(_00191_),
    .Q(\rvsingle.dp.rf.rf[18][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12734_ (.CLK(clknet_leaf_150_clk),
    .D(_00192_),
    .Q(\rvsingle.dp.rf.rf[18][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12735_ (.CLK(clknet_leaf_2_clk),
    .D(_00193_),
    .Q(\rvsingle.dp.rf.rf[18][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12736_ (.CLK(clknet_leaf_116_clk),
    .D(_00194_),
    .Q(\rvsingle.dp.rf.rf[18][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12737_ (.CLK(clknet_leaf_141_clk),
    .D(_00195_),
    .Q(\rvsingle.dp.rf.rf[18][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12738_ (.CLK(clknet_leaf_129_clk),
    .D(_00196_),
    .Q(\rvsingle.dp.rf.rf[18][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12739_ (.CLK(clknet_leaf_116_clk),
    .D(_00197_),
    .Q(\rvsingle.dp.rf.rf[18][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12740_ (.CLK(clknet_leaf_102_clk),
    .D(_00198_),
    .Q(\rvsingle.dp.rf.rf[18][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12741_ (.CLK(clknet_leaf_114_clk),
    .D(_00199_),
    .Q(\rvsingle.dp.rf.rf[18][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12742_ (.CLK(clknet_leaf_113_clk),
    .D(_00200_),
    .Q(\rvsingle.dp.rf.rf[18][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12743_ (.CLK(clknet_leaf_98_clk),
    .D(_00201_),
    .Q(\rvsingle.dp.rf.rf[18][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12744_ (.CLK(clknet_leaf_104_clk),
    .D(_00202_),
    .Q(\rvsingle.dp.rf.rf[18][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12745_ (.CLK(clknet_leaf_96_clk),
    .D(_00203_),
    .Q(\rvsingle.dp.rf.rf[18][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12746_ (.CLK(clknet_leaf_81_clk),
    .D(_00204_),
    .Q(\rvsingle.dp.rf.rf[18][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12747_ (.CLK(clknet_leaf_88_clk),
    .D(_00205_),
    .Q(\rvsingle.dp.rf.rf[31][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12748_ (.CLK(clknet_leaf_50_clk),
    .D(_00206_),
    .Q(\rvsingle.dp.rf.rf[31][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12749_ (.CLK(clknet_leaf_43_clk),
    .D(_00207_),
    .Q(\rvsingle.dp.rf.rf[31][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12750_ (.CLK(clknet_leaf_71_clk),
    .D(_00208_),
    .Q(\rvsingle.dp.rf.rf[31][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12751_ (.CLK(clknet_leaf_37_clk),
    .D(_00209_),
    .Q(\rvsingle.dp.rf.rf[31][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12752_ (.CLK(clknet_leaf_52_clk),
    .D(_00210_),
    .Q(\rvsingle.dp.rf.rf[31][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12753_ (.CLK(clknet_leaf_49_clk),
    .D(_00211_),
    .Q(\rvsingle.dp.rf.rf[31][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12754_ (.CLK(clknet_leaf_40_clk),
    .D(_00212_),
    .Q(\rvsingle.dp.rf.rf[31][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12755_ (.CLK(clknet_leaf_35_clk),
    .D(_00213_),
    .Q(\rvsingle.dp.rf.rf[31][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12756_ (.CLK(clknet_leaf_21_clk),
    .D(_00214_),
    .Q(\rvsingle.dp.rf.rf[31][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12757_ (.CLK(clknet_leaf_37_clk),
    .D(_00215_),
    .Q(\rvsingle.dp.rf.rf[31][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12758_ (.CLK(clknet_leaf_34_clk),
    .D(_00216_),
    .Q(\rvsingle.dp.rf.rf[31][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12759_ (.CLK(clknet_leaf_7_clk),
    .D(_00217_),
    .Q(\rvsingle.dp.rf.rf[31][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12760_ (.CLK(clknet_leaf_34_clk),
    .D(_00218_),
    .Q(\rvsingle.dp.rf.rf[31][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12761_ (.CLK(clknet_leaf_32_clk),
    .D(_00219_),
    .Q(\rvsingle.dp.rf.rf[31][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12762_ (.CLK(clknet_leaf_4_clk),
    .D(_00220_),
    .Q(\rvsingle.dp.rf.rf[31][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12763_ (.CLK(clknet_leaf_142_clk),
    .D(_00221_),
    .Q(\rvsingle.dp.rf.rf[31][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12764_ (.CLK(clknet_leaf_149_clk),
    .D(_00222_),
    .Q(\rvsingle.dp.rf.rf[31][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12765_ (.CLK(clknet_leaf_143_clk),
    .D(_00223_),
    .Q(\rvsingle.dp.rf.rf[31][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12766_ (.CLK(clknet_leaf_150_clk),
    .D(_00224_),
    .Q(\rvsingle.dp.rf.rf[31][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12767_ (.CLK(clknet_leaf_3_clk),
    .D(_00225_),
    .Q(\rvsingle.dp.rf.rf[31][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12768_ (.CLK(clknet_leaf_117_clk),
    .D(_00226_),
    .Q(\rvsingle.dp.rf.rf[31][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12769_ (.CLK(clknet_leaf_141_clk),
    .D(_00227_),
    .Q(\rvsingle.dp.rf.rf[31][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12770_ (.CLK(clknet_leaf_140_clk),
    .D(_00228_),
    .Q(\rvsingle.dp.rf.rf[31][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12771_ (.CLK(clknet_leaf_116_clk),
    .D(_00229_),
    .Q(\rvsingle.dp.rf.rf[31][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12772_ (.CLK(clknet_leaf_109_clk),
    .D(_00230_),
    .Q(\rvsingle.dp.rf.rf[31][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12773_ (.CLK(clknet_leaf_114_clk),
    .D(_00231_),
    .Q(\rvsingle.dp.rf.rf[31][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12774_ (.CLK(clknet_leaf_113_clk),
    .D(_00232_),
    .Q(\rvsingle.dp.rf.rf[31][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12775_ (.CLK(clknet_leaf_98_clk),
    .D(_00233_),
    .Q(\rvsingle.dp.rf.rf[31][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12776_ (.CLK(clknet_leaf_106_clk),
    .D(_00234_),
    .Q(\rvsingle.dp.rf.rf[31][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12777_ (.CLK(clknet_leaf_95_clk),
    .D(_00235_),
    .Q(\rvsingle.dp.rf.rf[31][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12778_ (.CLK(clknet_leaf_81_clk),
    .D(_00236_),
    .Q(\rvsingle.dp.rf.rf[31][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12779_ (.CLK(clknet_leaf_86_clk),
    .D(_00237_),
    .Q(\rvsingle.dp.rf.rf[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12780_ (.CLK(clknet_leaf_51_clk),
    .D(_00238_),
    .Q(\rvsingle.dp.rf.rf[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12781_ (.CLK(clknet_leaf_45_clk),
    .D(_00239_),
    .Q(\rvsingle.dp.rf.rf[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12782_ (.CLK(clknet_leaf_68_clk),
    .D(_00240_),
    .Q(\rvsingle.dp.rf.rf[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12783_ (.CLK(clknet_leaf_66_clk),
    .D(_00241_),
    .Q(\rvsingle.dp.rf.rf[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12784_ (.CLK(clknet_leaf_68_clk),
    .D(_00242_),
    .Q(\rvsingle.dp.rf.rf[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12785_ (.CLK(clknet_leaf_56_clk),
    .D(_00243_),
    .Q(\rvsingle.dp.rf.rf[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12786_ (.CLK(clknet_leaf_56_clk),
    .D(_00244_),
    .Q(\rvsingle.dp.rf.rf[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12787_ (.CLK(clknet_leaf_27_clk),
    .D(_00245_),
    .Q(\rvsingle.dp.rf.rf[17][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12788_ (.CLK(clknet_leaf_60_clk),
    .D(_00246_),
    .Q(\rvsingle.dp.rf.rf[17][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12789_ (.CLK(clknet_leaf_64_clk),
    .D(_00247_),
    .Q(\rvsingle.dp.rf.rf[17][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12790_ (.CLK(clknet_leaf_31_clk),
    .D(_00248_),
    .Q(\rvsingle.dp.rf.rf[17][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12791_ (.CLK(clknet_leaf_16_clk),
    .D(_00249_),
    .Q(\rvsingle.dp.rf.rf[17][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12792_ (.CLK(clknet_leaf_31_clk),
    .D(_00250_),
    .Q(\rvsingle.dp.rf.rf[17][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12793_ (.CLK(clknet_leaf_16_clk),
    .D(_00251_),
    .Q(\rvsingle.dp.rf.rf[17][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12794_ (.CLK(clknet_leaf_13_clk),
    .D(_00252_),
    .Q(\rvsingle.dp.rf.rf[17][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12795_ (.CLK(clknet_leaf_142_clk),
    .D(_00253_),
    .Q(\rvsingle.dp.rf.rf[17][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12796_ (.CLK(clknet_leaf_149_clk),
    .D(_00254_),
    .Q(\rvsingle.dp.rf.rf[17][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12797_ (.CLK(clknet_leaf_133_clk),
    .D(_00255_),
    .Q(\rvsingle.dp.rf.rf[17][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12798_ (.CLK(clknet_leaf_134_clk),
    .D(_00256_),
    .Q(\rvsingle.dp.rf.rf[17][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12799_ (.CLK(clknet_leaf_1_clk),
    .D(_00257_),
    .Q(\rvsingle.dp.rf.rf[17][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12800_ (.CLK(clknet_leaf_120_clk),
    .D(_00258_),
    .Q(\rvsingle.dp.rf.rf[17][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12801_ (.CLK(clknet_leaf_130_clk),
    .D(_00259_),
    .Q(\rvsingle.dp.rf.rf[17][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12802_ (.CLK(clknet_leaf_140_clk),
    .D(_00260_),
    .Q(\rvsingle.dp.rf.rf[17][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12803_ (.CLK(clknet_leaf_115_clk),
    .D(_00261_),
    .Q(\rvsingle.dp.rf.rf[17][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12804_ (.CLK(clknet_leaf_123_clk),
    .D(_00262_),
    .Q(\rvsingle.dp.rf.rf[17][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12805_ (.CLK(clknet_leaf_123_clk),
    .D(_00263_),
    .Q(\rvsingle.dp.rf.rf[17][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12806_ (.CLK(clknet_leaf_113_clk),
    .D(_00264_),
    .Q(\rvsingle.dp.rf.rf[17][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12807_ (.CLK(clknet_leaf_98_clk),
    .D(_00265_),
    .Q(\rvsingle.dp.rf.rf[17][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12808_ (.CLK(clknet_leaf_123_clk),
    .D(_00266_),
    .Q(\rvsingle.dp.rf.rf[17][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12809_ (.CLK(clknet_leaf_96_clk),
    .D(_00267_),
    .Q(\rvsingle.dp.rf.rf[17][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12810_ (.CLK(clknet_leaf_80_clk),
    .D(_00268_),
    .Q(\rvsingle.dp.rf.rf[17][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12811_ (.CLK(clknet_leaf_86_clk),
    .D(_00269_),
    .Q(\rvsingle.dp.rf.rf[16][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12812_ (.CLK(clknet_leaf_50_clk),
    .D(_00270_),
    .Q(\rvsingle.dp.rf.rf[16][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12813_ (.CLK(clknet_leaf_45_clk),
    .D(_00271_),
    .Q(\rvsingle.dp.rf.rf[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12814_ (.CLK(clknet_leaf_70_clk),
    .D(_00272_),
    .Q(\rvsingle.dp.rf.rf[16][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12815_ (.CLK(clknet_leaf_27_clk),
    .D(_00273_),
    .Q(\rvsingle.dp.rf.rf[16][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12816_ (.CLK(clknet_leaf_71_clk),
    .D(_00274_),
    .Q(\rvsingle.dp.rf.rf[16][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12817_ (.CLK(clknet_leaf_48_clk),
    .D(_00275_),
    .Q(\rvsingle.dp.rf.rf[16][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12818_ (.CLK(clknet_leaf_47_clk),
    .D(_00276_),
    .Q(\rvsingle.dp.rf.rf[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12819_ (.CLK(clknet_leaf_35_clk),
    .D(_00277_),
    .Q(\rvsingle.dp.rf.rf[16][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12820_ (.CLK(clknet_leaf_64_clk),
    .D(_00278_),
    .Q(\rvsingle.dp.rf.rf[16][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12821_ (.CLK(clknet_leaf_26_clk),
    .D(_00279_),
    .Q(\rvsingle.dp.rf.rf[16][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12822_ (.CLK(clknet_leaf_31_clk),
    .D(_00280_),
    .Q(\rvsingle.dp.rf.rf[16][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12823_ (.CLK(clknet_leaf_6_clk),
    .D(_00281_),
    .Q(\rvsingle.dp.rf.rf[16][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12824_ (.CLK(clknet_leaf_33_clk),
    .D(_00282_),
    .Q(\rvsingle.dp.rf.rf[16][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12825_ (.CLK(clknet_leaf_8_clk),
    .D(_00283_),
    .Q(\rvsingle.dp.rf.rf[16][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12826_ (.CLK(clknet_leaf_4_clk),
    .D(_00284_),
    .Q(\rvsingle.dp.rf.rf[16][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12827_ (.CLK(clknet_leaf_142_clk),
    .D(_00285_),
    .Q(\rvsingle.dp.rf.rf[16][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12828_ (.CLK(clknet_leaf_147_clk),
    .D(_00286_),
    .Q(\rvsingle.dp.rf.rf[16][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12829_ (.CLK(clknet_leaf_143_clk),
    .D(_00287_),
    .Q(\rvsingle.dp.rf.rf[16][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12830_ (.CLK(clknet_leaf_0_clk),
    .D(_00288_),
    .Q(\rvsingle.dp.rf.rf[16][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12831_ (.CLK(clknet_leaf_16_clk),
    .D(_00289_),
    .Q(\rvsingle.dp.rf.rf[16][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12832_ (.CLK(clknet_leaf_115_clk),
    .D(_00290_),
    .Q(\rvsingle.dp.rf.rf[16][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12833_ (.CLK(clknet_leaf_137_clk),
    .D(_00291_),
    .Q(\rvsingle.dp.rf.rf[16][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12834_ (.CLK(clknet_leaf_129_clk),
    .D(_00292_),
    .Q(\rvsingle.dp.rf.rf[16][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12835_ (.CLK(clknet_leaf_127_clk),
    .D(_00293_),
    .Q(\rvsingle.dp.rf.rf[16][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12836_ (.CLK(clknet_leaf_101_clk),
    .D(_00294_),
    .Q(\rvsingle.dp.rf.rf[16][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12837_ (.CLK(clknet_leaf_113_clk),
    .D(_00295_),
    .Q(\rvsingle.dp.rf.rf[16][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12838_ (.CLK(clknet_leaf_113_clk),
    .D(_00296_),
    .Q(\rvsingle.dp.rf.rf[16][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12839_ (.CLK(clknet_leaf_98_clk),
    .D(_00297_),
    .Q(\rvsingle.dp.rf.rf[16][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12840_ (.CLK(clknet_leaf_104_clk),
    .D(_00298_),
    .Q(\rvsingle.dp.rf.rf[16][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12841_ (.CLK(clknet_leaf_96_clk),
    .D(_00299_),
    .Q(\rvsingle.dp.rf.rf[16][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12842_ (.CLK(clknet_leaf_81_clk),
    .D(_00300_),
    .Q(\rvsingle.dp.rf.rf[16][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12843_ (.CLK(clknet_leaf_88_clk),
    .D(_00301_),
    .Q(\rvsingle.dp.rf.rf[29][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12844_ (.CLK(clknet_leaf_51_clk),
    .D(_00302_),
    .Q(\rvsingle.dp.rf.rf[29][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12845_ (.CLK(clknet_leaf_46_clk),
    .D(_00303_),
    .Q(\rvsingle.dp.rf.rf[29][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12846_ (.CLK(clknet_leaf_71_clk),
    .D(_00304_),
    .Q(\rvsingle.dp.rf.rf[29][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12847_ (.CLK(clknet_leaf_37_clk),
    .D(_00305_),
    .Q(\rvsingle.dp.rf.rf[29][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12848_ (.CLK(clknet_leaf_53_clk),
    .D(_00306_),
    .Q(\rvsingle.dp.rf.rf[29][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12849_ (.CLK(clknet_leaf_48_clk),
    .D(_00307_),
    .Q(\rvsingle.dp.rf.rf[29][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12850_ (.CLK(clknet_leaf_40_clk),
    .D(_00308_),
    .Q(\rvsingle.dp.rf.rf[29][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12851_ (.CLK(clknet_leaf_35_clk),
    .D(_00309_),
    .Q(\rvsingle.dp.rf.rf[29][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12852_ (.CLK(clknet_leaf_21_clk),
    .D(_00310_),
    .Q(\rvsingle.dp.rf.rf[29][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12853_ (.CLK(clknet_leaf_37_clk),
    .D(_00311_),
    .Q(\rvsingle.dp.rf.rf[29][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12854_ (.CLK(clknet_leaf_34_clk),
    .D(_00312_),
    .Q(\rvsingle.dp.rf.rf[29][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12855_ (.CLK(clknet_leaf_6_clk),
    .D(_00313_),
    .Q(\rvsingle.dp.rf.rf[29][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12856_ (.CLK(clknet_leaf_33_clk),
    .D(_00314_),
    .Q(\rvsingle.dp.rf.rf[29][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12857_ (.CLK(clknet_leaf_8_clk),
    .D(_00315_),
    .Q(\rvsingle.dp.rf.rf[29][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12858_ (.CLK(clknet_leaf_4_clk),
    .D(_00316_),
    .Q(\rvsingle.dp.rf.rf[29][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12859_ (.CLK(clknet_leaf_142_clk),
    .D(_00317_),
    .Q(\rvsingle.dp.rf.rf[29][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12860_ (.CLK(clknet_leaf_148_clk),
    .D(_00318_),
    .Q(\rvsingle.dp.rf.rf[29][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12861_ (.CLK(clknet_leaf_143_clk),
    .D(_00319_),
    .Q(\rvsingle.dp.rf.rf[29][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12862_ (.CLK(clknet_leaf_2_clk),
    .D(_00320_),
    .Q(\rvsingle.dp.rf.rf[29][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12863_ (.CLK(clknet_leaf_1_clk),
    .D(_00321_),
    .Q(\rvsingle.dp.rf.rf[29][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12864_ (.CLK(clknet_leaf_116_clk),
    .D(_00322_),
    .Q(\rvsingle.dp.rf.rf[29][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12865_ (.CLK(clknet_leaf_140_clk),
    .D(_00323_),
    .Q(\rvsingle.dp.rf.rf[29][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12866_ (.CLK(clknet_leaf_140_clk),
    .D(_00324_),
    .Q(\rvsingle.dp.rf.rf[29][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12867_ (.CLK(clknet_leaf_116_clk),
    .D(_00325_),
    .Q(\rvsingle.dp.rf.rf[29][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12868_ (.CLK(clknet_leaf_107_clk),
    .D(_00326_),
    .Q(\rvsingle.dp.rf.rf[29][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12869_ (.CLK(clknet_leaf_114_clk),
    .D(_00327_),
    .Q(\rvsingle.dp.rf.rf[29][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12870_ (.CLK(clknet_leaf_108_clk),
    .D(_00328_),
    .Q(\rvsingle.dp.rf.rf[29][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12871_ (.CLK(clknet_leaf_99_clk),
    .D(_00329_),
    .Q(\rvsingle.dp.rf.rf[29][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12872_ (.CLK(clknet_leaf_106_clk),
    .D(_00330_),
    .Q(\rvsingle.dp.rf.rf[29][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12873_ (.CLK(clknet_leaf_95_clk),
    .D(_00331_),
    .Q(\rvsingle.dp.rf.rf[29][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12874_ (.CLK(clknet_leaf_81_clk),
    .D(_00332_),
    .Q(\rvsingle.dp.rf.rf[29][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12875_ (.CLK(clknet_leaf_88_clk),
    .D(_00333_),
    .Q(\rvsingle.dp.rf.rf[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12876_ (.CLK(clknet_leaf_51_clk),
    .D(_00334_),
    .Q(\rvsingle.dp.rf.rf[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12877_ (.CLK(clknet_leaf_43_clk),
    .D(_00335_),
    .Q(\rvsingle.dp.rf.rf[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12878_ (.CLK(clknet_leaf_52_clk),
    .D(_00336_),
    .Q(\rvsingle.dp.rf.rf[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12879_ (.CLK(clknet_leaf_41_clk),
    .D(_00337_),
    .Q(\rvsingle.dp.rf.rf[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12880_ (.CLK(clknet_leaf_52_clk),
    .D(_00338_),
    .Q(\rvsingle.dp.rf.rf[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12881_ (.CLK(clknet_leaf_42_clk),
    .D(_00339_),
    .Q(\rvsingle.dp.rf.rf[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12882_ (.CLK(clknet_leaf_41_clk),
    .D(_00340_),
    .Q(\rvsingle.dp.rf.rf[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12883_ (.CLK(clknet_leaf_34_clk),
    .D(_00341_),
    .Q(\rvsingle.dp.rf.rf[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12884_ (.CLK(clknet_leaf_25_clk),
    .D(_00342_),
    .Q(\rvsingle.dp.rf.rf[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12885_ (.CLK(clknet_leaf_36_clk),
    .D(_00343_),
    .Q(\rvsingle.dp.rf.rf[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12886_ (.CLK(clknet_leaf_32_clk),
    .D(_00344_),
    .Q(\rvsingle.dp.rf.rf[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12887_ (.CLK(clknet_leaf_7_clk),
    .D(_00345_),
    .Q(\rvsingle.dp.rf.rf[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12888_ (.CLK(clknet_leaf_32_clk),
    .D(_00346_),
    .Q(\rvsingle.dp.rf.rf[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12889_ (.CLK(clknet_leaf_8_clk),
    .D(_00347_),
    .Q(\rvsingle.dp.rf.rf[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12890_ (.CLK(clknet_leaf_5_clk),
    .D(_00348_),
    .Q(\rvsingle.dp.rf.rf[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12891_ (.CLK(clknet_leaf_141_clk),
    .D(_00349_),
    .Q(\rvsingle.dp.rf.rf[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12892_ (.CLK(clknet_leaf_148_clk),
    .D(_00350_),
    .Q(\rvsingle.dp.rf.rf[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12893_ (.CLK(clknet_leaf_142_clk),
    .D(_00351_),
    .Q(\rvsingle.dp.rf.rf[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12894_ (.CLK(clknet_leaf_150_clk),
    .D(_00352_),
    .Q(\rvsingle.dp.rf.rf[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12895_ (.CLK(clknet_leaf_2_clk),
    .D(_00353_),
    .Q(\rvsingle.dp.rf.rf[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12896_ (.CLK(clknet_leaf_114_clk),
    .D(_00354_),
    .Q(\rvsingle.dp.rf.rf[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12897_ (.CLK(clknet_leaf_140_clk),
    .D(_00355_),
    .Q(\rvsingle.dp.rf.rf[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12898_ (.CLK(clknet_leaf_141_clk),
    .D(_00356_),
    .Q(\rvsingle.dp.rf.rf[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12899_ (.CLK(clknet_leaf_116_clk),
    .D(_00357_),
    .Q(\rvsingle.dp.rf.rf[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12900_ (.CLK(clknet_leaf_110_clk),
    .D(_00358_),
    .Q(\rvsingle.dp.rf.rf[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12901_ (.CLK(clknet_leaf_108_clk),
    .D(_00359_),
    .Q(\rvsingle.dp.rf.rf[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12902_ (.CLK(clknet_leaf_114_clk),
    .D(_00360_),
    .Q(\rvsingle.dp.rf.rf[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12903_ (.CLK(clknet_leaf_98_clk),
    .D(_00361_),
    .Q(\rvsingle.dp.rf.rf[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12904_ (.CLK(clknet_leaf_105_clk),
    .D(_00362_),
    .Q(\rvsingle.dp.rf.rf[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12905_ (.CLK(clknet_leaf_97_clk),
    .D(_00363_),
    .Q(\rvsingle.dp.rf.rf[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12906_ (.CLK(clknet_leaf_95_clk),
    .D(_00364_),
    .Q(\rvsingle.dp.rf.rf[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12907_ (.CLK(clknet_leaf_88_clk),
    .D(_00365_),
    .Q(\rvsingle.dp.rf.rf[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12908_ (.CLK(clknet_leaf_50_clk),
    .D(_00366_),
    .Q(\rvsingle.dp.rf.rf[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12909_ (.CLK(clknet_leaf_43_clk),
    .D(_00367_),
    .Q(\rvsingle.dp.rf.rf[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12910_ (.CLK(clknet_leaf_52_clk),
    .D(_00368_),
    .Q(\rvsingle.dp.rf.rf[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12911_ (.CLK(clknet_leaf_40_clk),
    .D(_00369_),
    .Q(\rvsingle.dp.rf.rf[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12912_ (.CLK(clknet_leaf_52_clk),
    .D(_00370_),
    .Q(\rvsingle.dp.rf.rf[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12913_ (.CLK(clknet_leaf_42_clk),
    .D(_00371_),
    .Q(\rvsingle.dp.rf.rf[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12914_ (.CLK(clknet_leaf_40_clk),
    .D(_00372_),
    .Q(\rvsingle.dp.rf.rf[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12915_ (.CLK(clknet_leaf_34_clk),
    .D(_00373_),
    .Q(\rvsingle.dp.rf.rf[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12916_ (.CLK(clknet_leaf_61_clk),
    .D(_00374_),
    .Q(\rvsingle.dp.rf.rf[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12917_ (.CLK(clknet_leaf_37_clk),
    .D(_00375_),
    .Q(\rvsingle.dp.rf.rf[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12918_ (.CLK(clknet_leaf_32_clk),
    .D(_00376_),
    .Q(\rvsingle.dp.rf.rf[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12919_ (.CLK(clknet_leaf_7_clk),
    .D(_00377_),
    .Q(\rvsingle.dp.rf.rf[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12920_ (.CLK(clknet_leaf_32_clk),
    .D(_00378_),
    .Q(\rvsingle.dp.rf.rf[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12921_ (.CLK(clknet_leaf_8_clk),
    .D(_00379_),
    .Q(\rvsingle.dp.rf.rf[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12922_ (.CLK(clknet_leaf_3_clk),
    .D(_00380_),
    .Q(\rvsingle.dp.rf.rf[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12923_ (.CLK(clknet_leaf_141_clk),
    .D(_00381_),
    .Q(\rvsingle.dp.rf.rf[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12924_ (.CLK(clknet_leaf_148_clk),
    .D(_00382_),
    .Q(\rvsingle.dp.rf.rf[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12925_ (.CLK(clknet_leaf_142_clk),
    .D(_00383_),
    .Q(\rvsingle.dp.rf.rf[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12926_ (.CLK(clknet_leaf_150_clk),
    .D(_00384_),
    .Q(\rvsingle.dp.rf.rf[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12927_ (.CLK(clknet_leaf_2_clk),
    .D(_00385_),
    .Q(\rvsingle.dp.rf.rf[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12928_ (.CLK(clknet_leaf_116_clk),
    .D(_00386_),
    .Q(\rvsingle.dp.rf.rf[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12929_ (.CLK(clknet_leaf_117_clk),
    .D(_00387_),
    .Q(\rvsingle.dp.rf.rf[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12930_ (.CLK(clknet_leaf_141_clk),
    .D(_00388_),
    .Q(\rvsingle.dp.rf.rf[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12931_ (.CLK(clknet_leaf_116_clk),
    .D(_00389_),
    .Q(\rvsingle.dp.rf.rf[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12932_ (.CLK(clknet_leaf_110_clk),
    .D(_00390_),
    .Q(\rvsingle.dp.rf.rf[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12933_ (.CLK(clknet_leaf_108_clk),
    .D(_00391_),
    .Q(\rvsingle.dp.rf.rf[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12934_ (.CLK(clknet_leaf_114_clk),
    .D(_00392_),
    .Q(\rvsingle.dp.rf.rf[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12935_ (.CLK(clknet_leaf_98_clk),
    .D(_00393_),
    .Q(\rvsingle.dp.rf.rf[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12936_ (.CLK(clknet_leaf_105_clk),
    .D(_00394_),
    .Q(\rvsingle.dp.rf.rf[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12937_ (.CLK(clknet_leaf_97_clk),
    .D(_00395_),
    .Q(\rvsingle.dp.rf.rf[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12938_ (.CLK(clknet_leaf_81_clk),
    .D(_00396_),
    .Q(\rvsingle.dp.rf.rf[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12939_ (.CLK(clknet_leaf_86_clk),
    .D(_00397_),
    .Q(\rvsingle.dp.rf.rf[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12940_ (.CLK(clknet_leaf_52_clk),
    .D(_00398_),
    .Q(\rvsingle.dp.rf.rf[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12941_ (.CLK(clknet_leaf_42_clk),
    .D(_00399_),
    .Q(\rvsingle.dp.rf.rf[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12942_ (.CLK(clknet_leaf_52_clk),
    .D(_00400_),
    .Q(\rvsingle.dp.rf.rf[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12943_ (.CLK(clknet_leaf_40_clk),
    .D(_00401_),
    .Q(\rvsingle.dp.rf.rf[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12944_ (.CLK(clknet_leaf_51_clk),
    .D(_00402_),
    .Q(\rvsingle.dp.rf.rf[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12945_ (.CLK(clknet_leaf_42_clk),
    .D(_00403_),
    .Q(\rvsingle.dp.rf.rf[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12946_ (.CLK(clknet_leaf_41_clk),
    .D(_00404_),
    .Q(\rvsingle.dp.rf.rf[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12947_ (.CLK(clknet_leaf_34_clk),
    .D(_00405_),
    .Q(\rvsingle.dp.rf.rf[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12948_ (.CLK(clknet_leaf_22_clk),
    .D(_00406_),
    .Q(\rvsingle.dp.rf.rf[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12949_ (.CLK(clknet_leaf_36_clk),
    .D(_00407_),
    .Q(\rvsingle.dp.rf.rf[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12950_ (.CLK(clknet_leaf_31_clk),
    .D(_00408_),
    .Q(\rvsingle.dp.rf.rf[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12951_ (.CLK(clknet_leaf_9_clk),
    .D(_00409_),
    .Q(\rvsingle.dp.rf.rf[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12952_ (.CLK(clknet_leaf_23_clk),
    .D(_00410_),
    .Q(\rvsingle.dp.rf.rf[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12953_ (.CLK(clknet_leaf_9_clk),
    .D(_00411_),
    .Q(\rvsingle.dp.rf.rf[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12954_ (.CLK(clknet_leaf_1_clk),
    .D(_00412_),
    .Q(\rvsingle.dp.rf.rf[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12955_ (.CLK(clknet_leaf_141_clk),
    .D(_00413_),
    .Q(\rvsingle.dp.rf.rf[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12956_ (.CLK(clknet_leaf_148_clk),
    .D(_00414_),
    .Q(\rvsingle.dp.rf.rf[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12957_ (.CLK(clknet_leaf_142_clk),
    .D(_00415_),
    .Q(\rvsingle.dp.rf.rf[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12958_ (.CLK(clknet_leaf_150_clk),
    .D(_00416_),
    .Q(\rvsingle.dp.rf.rf[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12959_ (.CLK(clknet_leaf_2_clk),
    .D(_00417_),
    .Q(\rvsingle.dp.rf.rf[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12960_ (.CLK(clknet_leaf_115_clk),
    .D(_00418_),
    .Q(\rvsingle.dp.rf.rf[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12961_ (.CLK(clknet_leaf_140_clk),
    .D(_00419_),
    .Q(\rvsingle.dp.rf.rf[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12962_ (.CLK(clknet_leaf_141_clk),
    .D(_00420_),
    .Q(\rvsingle.dp.rf.rf[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12963_ (.CLK(clknet_leaf_116_clk),
    .D(_00421_),
    .Q(\rvsingle.dp.rf.rf[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12964_ (.CLK(clknet_leaf_110_clk),
    .D(_00422_),
    .Q(\rvsingle.dp.rf.rf[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12965_ (.CLK(clknet_leaf_108_clk),
    .D(_00423_),
    .Q(\rvsingle.dp.rf.rf[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12966_ (.CLK(clknet_leaf_114_clk),
    .D(_00424_),
    .Q(\rvsingle.dp.rf.rf[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12967_ (.CLK(clknet_leaf_98_clk),
    .D(_00425_),
    .Q(\rvsingle.dp.rf.rf[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 _12968_ (.CLK(clknet_leaf_105_clk),
    .D(_00426_),
    .Q(\rvsingle.dp.rf.rf[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 _12969_ (.CLK(clknet_leaf_97_clk),
    .D(_00427_),
    .Q(\rvsingle.dp.rf.rf[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _12970_ (.CLK(clknet_leaf_81_clk),
    .D(_00428_),
    .Q(\rvsingle.dp.rf.rf[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _12971_ (.CLK(clknet_leaf_86_clk),
    .D(_00429_),
    .Q(\rvsingle.dp.rf.rf[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _12972_ (.CLK(clknet_leaf_52_clk),
    .D(_00430_),
    .Q(\rvsingle.dp.rf.rf[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _12973_ (.CLK(clknet_leaf_42_clk),
    .D(_00431_),
    .Q(\rvsingle.dp.rf.rf[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _12974_ (.CLK(clknet_leaf_52_clk),
    .D(_00432_),
    .Q(\rvsingle.dp.rf.rf[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _12975_ (.CLK(clknet_leaf_40_clk),
    .D(_00433_),
    .Q(\rvsingle.dp.rf.rf[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _12976_ (.CLK(clknet_leaf_52_clk),
    .D(_00434_),
    .Q(\rvsingle.dp.rf.rf[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _12977_ (.CLK(clknet_leaf_40_clk),
    .D(_00435_),
    .Q(\rvsingle.dp.rf.rf[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _12978_ (.CLK(clknet_leaf_40_clk),
    .D(_00436_),
    .Q(\rvsingle.dp.rf.rf[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _12979_ (.CLK(clknet_leaf_34_clk),
    .D(_00437_),
    .Q(\rvsingle.dp.rf.rf[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _12980_ (.CLK(clknet_leaf_22_clk),
    .D(_00438_),
    .Q(\rvsingle.dp.rf.rf[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _12981_ (.CLK(clknet_leaf_37_clk),
    .D(_00439_),
    .Q(\rvsingle.dp.rf.rf[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _12982_ (.CLK(clknet_leaf_31_clk),
    .D(_00440_),
    .Q(\rvsingle.dp.rf.rf[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _12983_ (.CLK(clknet_leaf_9_clk),
    .D(_00441_),
    .Q(\rvsingle.dp.rf.rf[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _12984_ (.CLK(clknet_leaf_23_clk),
    .D(_00442_),
    .Q(\rvsingle.dp.rf.rf[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _12985_ (.CLK(clknet_leaf_9_clk),
    .D(_00443_),
    .Q(\rvsingle.dp.rf.rf[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _12986_ (.CLK(clknet_leaf_1_clk),
    .D(_00444_),
    .Q(\rvsingle.dp.rf.rf[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _12987_ (.CLK(clknet_leaf_141_clk),
    .D(_00445_),
    .Q(\rvsingle.dp.rf.rf[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _12988_ (.CLK(clknet_leaf_148_clk),
    .D(_00446_),
    .Q(\rvsingle.dp.rf.rf[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _12989_ (.CLK(clknet_leaf_142_clk),
    .D(_00447_),
    .Q(\rvsingle.dp.rf.rf[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _12990_ (.CLK(clknet_leaf_150_clk),
    .D(_00448_),
    .Q(\rvsingle.dp.rf.rf[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _12991_ (.CLK(clknet_leaf_2_clk),
    .D(_00449_),
    .Q(\rvsingle.dp.rf.rf[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _12992_ (.CLK(clknet_leaf_115_clk),
    .D(_00450_),
    .Q(\rvsingle.dp.rf.rf[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _12993_ (.CLK(clknet_leaf_140_clk),
    .D(_00451_),
    .Q(\rvsingle.dp.rf.rf[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _12994_ (.CLK(clknet_leaf_141_clk),
    .D(_00452_),
    .Q(\rvsingle.dp.rf.rf[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _12995_ (.CLK(clknet_leaf_116_clk),
    .D(_00453_),
    .Q(\rvsingle.dp.rf.rf[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _12996_ (.CLK(clknet_leaf_109_clk),
    .D(_00454_),
    .Q(\rvsingle.dp.rf.rf[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _12997_ (.CLK(clknet_leaf_108_clk),
    .D(_00455_),
    .Q(\rvsingle.dp.rf.rf[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 _12998_ (.CLK(clknet_leaf_115_clk),
    .D(_00456_),
    .Q(\rvsingle.dp.rf.rf[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _12999_ (.CLK(clknet_leaf_98_clk),
    .D(_00457_),
    .Q(\rvsingle.dp.rf.rf[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13000_ (.CLK(clknet_leaf_105_clk),
    .D(_00458_),
    .Q(\rvsingle.dp.rf.rf[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13001_ (.CLK(clknet_leaf_97_clk),
    .D(_00459_),
    .Q(\rvsingle.dp.rf.rf[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13002_ (.CLK(clknet_leaf_81_clk),
    .D(_00460_),
    .Q(\rvsingle.dp.rf.rf[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13003_ (.CLK(clknet_leaf_89_clk),
    .D(_00461_),
    .Q(\rvsingle.dp.rf.rf[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13004_ (.CLK(clknet_leaf_51_clk),
    .D(_00462_),
    .Q(\rvsingle.dp.rf.rf[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13005_ (.CLK(clknet_leaf_45_clk),
    .D(_00463_),
    .Q(\rvsingle.dp.rf.rf[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13006_ (.CLK(clknet_leaf_55_clk),
    .D(_00464_),
    .Q(\rvsingle.dp.rf.rf[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13007_ (.CLK(clknet_leaf_57_clk),
    .D(_00465_),
    .Q(\rvsingle.dp.rf.rf[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13008_ (.CLK(clknet_leaf_55_clk),
    .D(_00466_),
    .Q(\rvsingle.dp.rf.rf[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13009_ (.CLK(clknet_leaf_57_clk),
    .D(_00467_),
    .Q(\rvsingle.dp.rf.rf[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13010_ (.CLK(clknet_leaf_57_clk),
    .D(_00468_),
    .Q(\rvsingle.dp.rf.rf[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13011_ (.CLK(clknet_leaf_29_clk),
    .D(_00469_),
    .Q(\rvsingle.dp.rf.rf[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13012_ (.CLK(clknet_leaf_61_clk),
    .D(_00470_),
    .Q(\rvsingle.dp.rf.rf[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13013_ (.CLK(clknet_leaf_65_clk),
    .D(_00471_),
    .Q(\rvsingle.dp.rf.rf[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13014_ (.CLK(clknet_leaf_25_clk),
    .D(_00472_),
    .Q(\rvsingle.dp.rf.rf[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13015_ (.CLK(clknet_leaf_11_clk),
    .D(_00473_),
    .Q(\rvsingle.dp.rf.rf[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13016_ (.CLK(clknet_leaf_23_clk),
    .D(_00474_),
    .Q(\rvsingle.dp.rf.rf[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13017_ (.CLK(clknet_leaf_10_clk),
    .D(_00475_),
    .Q(\rvsingle.dp.rf.rf[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13018_ (.CLK(clknet_leaf_12_clk),
    .D(_00476_),
    .Q(\rvsingle.dp.rf.rf[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13019_ (.CLK(clknet_leaf_136_clk),
    .D(_00477_),
    .Q(\rvsingle.dp.rf.rf[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13020_ (.CLK(clknet_leaf_13_clk),
    .D(_00478_),
    .Q(\rvsingle.dp.rf.rf[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13021_ (.CLK(clknet_leaf_145_clk),
    .D(_00479_),
    .Q(\rvsingle.dp.rf.rf[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13022_ (.CLK(clknet_leaf_134_clk),
    .D(_00480_),
    .Q(\rvsingle.dp.rf.rf[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13023_ (.CLK(clknet_leaf_13_clk),
    .D(_00481_),
    .Q(\rvsingle.dp.rf.rf[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13024_ (.CLK(clknet_leaf_118_clk),
    .D(_00482_),
    .Q(\rvsingle.dp.rf.rf[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13025_ (.CLK(clknet_leaf_126_clk),
    .D(_00483_),
    .Q(\rvsingle.dp.rf.rf[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13026_ (.CLK(clknet_leaf_132_clk),
    .D(_00484_),
    .Q(\rvsingle.dp.rf.rf[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13027_ (.CLK(clknet_leaf_125_clk),
    .D(_00485_),
    .Q(\rvsingle.dp.rf.rf[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13028_ (.CLK(clknet_leaf_124_clk),
    .D(_00486_),
    .Q(\rvsingle.dp.rf.rf[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13029_ (.CLK(clknet_leaf_111_clk),
    .D(_00487_),
    .Q(\rvsingle.dp.rf.rf[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13030_ (.CLK(clknet_leaf_112_clk),
    .D(_00488_),
    .Q(\rvsingle.dp.rf.rf[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13031_ (.CLK(clknet_leaf_101_clk),
    .D(_00489_),
    .Q(\rvsingle.dp.rf.rf[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13032_ (.CLK(clknet_leaf_102_clk),
    .D(_00490_),
    .Q(\rvsingle.dp.rf.rf[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13033_ (.CLK(clknet_leaf_90_clk),
    .D(_00491_),
    .Q(\rvsingle.dp.rf.rf[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13034_ (.CLK(clknet_leaf_93_clk),
    .D(_00492_),
    .Q(\rvsingle.dp.rf.rf[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13035_ (.CLK(clknet_leaf_87_clk),
    .D(_00493_),
    .Q(\rvsingle.dp.rf.rf[19][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13036_ (.CLK(clknet_leaf_50_clk),
    .D(_00494_),
    .Q(\rvsingle.dp.rf.rf[19][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13037_ (.CLK(clknet_leaf_44_clk),
    .D(_00495_),
    .Q(\rvsingle.dp.rf.rf[19][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13038_ (.CLK(clknet_4_15_0_clk),
    .D(_00496_),
    .Q(\rvsingle.dp.rf.rf[19][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13039_ (.CLK(clknet_leaf_57_clk),
    .D(_00497_),
    .Q(\rvsingle.dp.rf.rf[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13040_ (.CLK(clknet_leaf_55_clk),
    .D(_00498_),
    .Q(\rvsingle.dp.rf.rf[19][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13041_ (.CLK(clknet_leaf_57_clk),
    .D(_00499_),
    .Q(\rvsingle.dp.rf.rf[19][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13042_ (.CLK(clknet_leaf_57_clk),
    .D(_00500_),
    .Q(\rvsingle.dp.rf.rf[19][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13043_ (.CLK(clknet_leaf_26_clk),
    .D(_00501_),
    .Q(\rvsingle.dp.rf.rf[19][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13044_ (.CLK(clknet_leaf_61_clk),
    .D(_00502_),
    .Q(\rvsingle.dp.rf.rf[19][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13045_ (.CLK(clknet_leaf_58_clk),
    .D(_00503_),
    .Q(\rvsingle.dp.rf.rf[19][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13046_ (.CLK(clknet_leaf_23_clk),
    .D(_00504_),
    .Q(\rvsingle.dp.rf.rf[19][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13047_ (.CLK(clknet_leaf_11_clk),
    .D(_00505_),
    .Q(\rvsingle.dp.rf.rf[19][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13048_ (.CLK(clknet_leaf_10_clk),
    .D(_00506_),
    .Q(\rvsingle.dp.rf.rf[19][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13049_ (.CLK(clknet_leaf_10_clk),
    .D(_00507_),
    .Q(\rvsingle.dp.rf.rf[19][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13050_ (.CLK(clknet_leaf_12_clk),
    .D(_00508_),
    .Q(\rvsingle.dp.rf.rf[19][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13051_ (.CLK(clknet_leaf_131_clk),
    .D(_00509_),
    .Q(\rvsingle.dp.rf.rf[19][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13052_ (.CLK(clknet_leaf_13_clk),
    .D(_00510_),
    .Q(\rvsingle.dp.rf.rf[19][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13053_ (.CLK(clknet_leaf_143_clk),
    .D(_00511_),
    .Q(\rvsingle.dp.rf.rf[19][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13054_ (.CLK(clknet_leaf_134_clk),
    .D(_00512_),
    .Q(\rvsingle.dp.rf.rf[19][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13055_ (.CLK(clknet_leaf_13_clk),
    .D(_00513_),
    .Q(\rvsingle.dp.rf.rf[19][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13056_ (.CLK(clknet_leaf_116_clk),
    .D(_00514_),
    .Q(\rvsingle.dp.rf.rf[19][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13057_ (.CLK(clknet_leaf_126_clk),
    .D(_00515_),
    .Q(\rvsingle.dp.rf.rf[19][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13058_ (.CLK(clknet_leaf_129_clk),
    .D(_00516_),
    .Q(\rvsingle.dp.rf.rf[19][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13059_ (.CLK(clknet_leaf_125_clk),
    .D(_00517_),
    .Q(\rvsingle.dp.rf.rf[19][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13060_ (.CLK(clknet_leaf_123_clk),
    .D(_00518_),
    .Q(\rvsingle.dp.rf.rf[19][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13061_ (.CLK(clknet_leaf_114_clk),
    .D(_00519_),
    .Q(\rvsingle.dp.rf.rf[19][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13062_ (.CLK(clknet_leaf_113_clk),
    .D(_00520_),
    .Q(\rvsingle.dp.rf.rf[19][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13063_ (.CLK(clknet_leaf_97_clk),
    .D(_00521_),
    .Q(\rvsingle.dp.rf.rf[19][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13064_ (.CLK(clknet_leaf_103_clk),
    .D(_00522_),
    .Q(\rvsingle.dp.rf.rf[19][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13065_ (.CLK(clknet_leaf_89_clk),
    .D(_00523_),
    .Q(\rvsingle.dp.rf.rf[19][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13066_ (.CLK(clknet_leaf_82_clk),
    .D(_00524_),
    .Q(\rvsingle.dp.rf.rf[19][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13067_ (.CLK(clknet_leaf_90_clk),
    .D(_00525_),
    .Q(\rvsingle.dp.rf.rf[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13068_ (.CLK(clknet_leaf_51_clk),
    .D(_00526_),
    .Q(\rvsingle.dp.rf.rf[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13069_ (.CLK(clknet_leaf_43_clk),
    .D(_00527_),
    .Q(\rvsingle.dp.rf.rf[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13070_ (.CLK(clknet_leaf_52_clk),
    .D(_00528_),
    .Q(\rvsingle.dp.rf.rf[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13071_ (.CLK(clknet_leaf_27_clk),
    .D(_00529_),
    .Q(\rvsingle.dp.rf.rf[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13072_ (.CLK(clknet_leaf_51_clk),
    .D(_00530_),
    .Q(\rvsingle.dp.rf.rf[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13073_ (.CLK(clknet_leaf_48_clk),
    .D(_00531_),
    .Q(\rvsingle.dp.rf.rf[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13074_ (.CLK(clknet_leaf_57_clk),
    .D(_00532_),
    .Q(\rvsingle.dp.rf.rf[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13075_ (.CLK(clknet_leaf_29_clk),
    .D(_00533_),
    .Q(\rvsingle.dp.rf.rf[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13076_ (.CLK(clknet_leaf_21_clk),
    .D(_00534_),
    .Q(\rvsingle.dp.rf.rf[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13077_ (.CLK(clknet_leaf_65_clk),
    .D(_00535_),
    .Q(\rvsingle.dp.rf.rf[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13078_ (.CLK(clknet_leaf_24_clk),
    .D(_00536_),
    .Q(\rvsingle.dp.rf.rf[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13079_ (.CLK(clknet_leaf_10_clk),
    .D(_00537_),
    .Q(\rvsingle.dp.rf.rf[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13080_ (.CLK(clknet_leaf_22_clk),
    .D(_00538_),
    .Q(\rvsingle.dp.rf.rf[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13081_ (.CLK(clknet_leaf_9_clk),
    .D(_00539_),
    .Q(\rvsingle.dp.rf.rf[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13082_ (.CLK(clknet_leaf_6_clk),
    .D(_00540_),
    .Q(\rvsingle.dp.rf.rf[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13083_ (.CLK(clknet_leaf_135_clk),
    .D(_00541_),
    .Q(\rvsingle.dp.rf.rf[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13084_ (.CLK(clknet_leaf_151_clk),
    .D(_00542_),
    .Q(\rvsingle.dp.rf.rf[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13085_ (.CLK(clknet_leaf_146_clk),
    .D(_00543_),
    .Q(\rvsingle.dp.rf.rf[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13086_ (.CLK(clknet_leaf_0_clk),
    .D(_00544_),
    .Q(\rvsingle.dp.rf.rf[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13087_ (.CLK(clknet_leaf_2_clk),
    .D(_00545_),
    .Q(\rvsingle.dp.rf.rf[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13088_ (.CLK(clknet_leaf_119_clk),
    .D(_00546_),
    .Q(\rvsingle.dp.rf.rf[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13089_ (.CLK(clknet_leaf_137_clk),
    .D(_00547_),
    .Q(\rvsingle.dp.rf.rf[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13090_ (.CLK(clknet_leaf_129_clk),
    .D(_00548_),
    .Q(\rvsingle.dp.rf.rf[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13091_ (.CLK(clknet_leaf_120_clk),
    .D(_00549_),
    .Q(\rvsingle.dp.rf.rf[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13092_ (.CLK(clknet_leaf_101_clk),
    .D(_00550_),
    .Q(\rvsingle.dp.rf.rf[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13093_ (.CLK(clknet_leaf_110_clk),
    .D(_00551_),
    .Q(\rvsingle.dp.rf.rf[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13094_ (.CLK(clknet_leaf_121_clk),
    .D(_00552_),
    .Q(\rvsingle.dp.rf.rf[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13095_ (.CLK(clknet_leaf_101_clk),
    .D(_00553_),
    .Q(\rvsingle.dp.rf.rf[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13096_ (.CLK(clknet_leaf_102_clk),
    .D(_00554_),
    .Q(\rvsingle.dp.rf.rf[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13097_ (.CLK(clknet_leaf_92_clk),
    .D(_00555_),
    .Q(\rvsingle.dp.rf.rf[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13098_ (.CLK(clknet_leaf_82_clk),
    .D(_00556_),
    .Q(\rvsingle.dp.rf.rf[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13099_ (.CLK(clknet_leaf_88_clk),
    .D(_00557_),
    .Q(\rvsingle.dp.rf.rf[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13100_ (.CLK(clknet_leaf_53_clk),
    .D(_00558_),
    .Q(\rvsingle.dp.rf.rf[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13101_ (.CLK(clknet_leaf_44_clk),
    .D(_00559_),
    .Q(\rvsingle.dp.rf.rf[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13102_ (.CLK(clknet_leaf_55_clk),
    .D(_00560_),
    .Q(\rvsingle.dp.rf.rf[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13103_ (.CLK(clknet_leaf_58_clk),
    .D(_00561_),
    .Q(\rvsingle.dp.rf.rf[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13104_ (.CLK(clknet_leaf_51_clk),
    .D(_00562_),
    .Q(\rvsingle.dp.rf.rf[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13105_ (.CLK(clknet_leaf_57_clk),
    .D(_00563_),
    .Q(\rvsingle.dp.rf.rf[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13106_ (.CLK(clknet_leaf_56_clk),
    .D(_00564_),
    .Q(\rvsingle.dp.rf.rf[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13107_ (.CLK(clknet_leaf_16_clk),
    .D(_00565_),
    .Q(\rvsingle.dp.rf.rf[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13108_ (.CLK(clknet_leaf_61_clk),
    .D(_00566_),
    .Q(\rvsingle.dp.rf.rf[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13109_ (.CLK(clknet_leaf_65_clk),
    .D(_00567_),
    .Q(\rvsingle.dp.rf.rf[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13110_ (.CLK(clknet_leaf_25_clk),
    .D(_00568_),
    .Q(\rvsingle.dp.rf.rf[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13111_ (.CLK(clknet_leaf_15_clk),
    .D(_00569_),
    .Q(\rvsingle.dp.rf.rf[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13112_ (.CLK(clknet_leaf_18_clk),
    .D(_00570_),
    .Q(\rvsingle.dp.rf.rf[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13113_ (.CLK(clknet_leaf_18_clk),
    .D(_00571_),
    .Q(\rvsingle.dp.rf.rf[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13114_ (.CLK(clknet_leaf_14_clk),
    .D(_00572_),
    .Q(\rvsingle.dp.rf.rf[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13115_ (.CLK(clknet_leaf_131_clk),
    .D(_00573_),
    .Q(\rvsingle.dp.rf.rf[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13116_ (.CLK(clknet_leaf_13_clk),
    .D(_00574_),
    .Q(\rvsingle.dp.rf.rf[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13117_ (.CLK(clknet_leaf_145_clk),
    .D(_00575_),
    .Q(\rvsingle.dp.rf.rf[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13118_ (.CLK(clknet_leaf_133_clk),
    .D(_00576_),
    .Q(\rvsingle.dp.rf.rf[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13119_ (.CLK(clknet_leaf_133_clk),
    .D(_00577_),
    .Q(\rvsingle.dp.rf.rf[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13120_ (.CLK(clknet_leaf_138_clk),
    .D(_00578_),
    .Q(\rvsingle.dp.rf.rf[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13121_ (.CLK(clknet_leaf_126_clk),
    .D(_00579_),
    .Q(\rvsingle.dp.rf.rf[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13122_ (.CLK(clknet_leaf_136_clk),
    .D(_00580_),
    .Q(\rvsingle.dp.rf.rf[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13123_ (.CLK(clknet_leaf_123_clk),
    .D(_00581_),
    .Q(\rvsingle.dp.rf.rf[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13124_ (.CLK(clknet_leaf_124_clk),
    .D(_00582_),
    .Q(\rvsingle.dp.rf.rf[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13125_ (.CLK(clknet_leaf_101_clk),
    .D(_00583_),
    .Q(\rvsingle.dp.rf.rf[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13126_ (.CLK(clknet_leaf_111_clk),
    .D(_00584_),
    .Q(\rvsingle.dp.rf.rf[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13127_ (.CLK(clknet_leaf_92_clk),
    .D(_00585_),
    .Q(\rvsingle.dp.rf.rf[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13128_ (.CLK(clknet_leaf_101_clk),
    .D(_00586_),
    .Q(\rvsingle.dp.rf.rf[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13129_ (.CLK(clknet_leaf_92_clk),
    .D(_00587_),
    .Q(\rvsingle.dp.rf.rf[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13130_ (.CLK(clknet_leaf_93_clk),
    .D(_00588_),
    .Q(\rvsingle.dp.rf.rf[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13131_ (.CLK(clknet_leaf_87_clk),
    .D(_00589_),
    .Q(\rvsingle.dp.rf.rf[23][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13132_ (.CLK(clknet_leaf_48_clk),
    .D(_00590_),
    .Q(\rvsingle.dp.rf.rf[23][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13133_ (.CLK(clknet_leaf_45_clk),
    .D(_00591_),
    .Q(\rvsingle.dp.rf.rf[23][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13134_ (.CLK(clknet_leaf_71_clk),
    .D(_00592_),
    .Q(\rvsingle.dp.rf.rf[23][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13135_ (.CLK(clknet_leaf_37_clk),
    .D(_00593_),
    .Q(\rvsingle.dp.rf.rf[23][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13136_ (.CLK(clknet_leaf_71_clk),
    .D(_00594_),
    .Q(\rvsingle.dp.rf.rf[23][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13137_ (.CLK(clknet_leaf_48_clk),
    .D(_00595_),
    .Q(\rvsingle.dp.rf.rf[23][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13138_ (.CLK(clknet_leaf_40_clk),
    .D(_00596_),
    .Q(\rvsingle.dp.rf.rf[23][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13139_ (.CLK(clknet_leaf_28_clk),
    .D(_00597_),
    .Q(\rvsingle.dp.rf.rf[23][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13140_ (.CLK(clknet_leaf_58_clk),
    .D(_00598_),
    .Q(\rvsingle.dp.rf.rf[23][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13141_ (.CLK(clknet_leaf_37_clk),
    .D(_00599_),
    .Q(\rvsingle.dp.rf.rf[23][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13142_ (.CLK(clknet_leaf_31_clk),
    .D(_00600_),
    .Q(\rvsingle.dp.rf.rf[23][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13143_ (.CLK(clknet_leaf_9_clk),
    .D(_00601_),
    .Q(\rvsingle.dp.rf.rf[23][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13144_ (.CLK(clknet_leaf_28_clk),
    .D(_00602_),
    .Q(\rvsingle.dp.rf.rf[23][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13145_ (.CLK(clknet_leaf_9_clk),
    .D(_00603_),
    .Q(\rvsingle.dp.rf.rf[23][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13146_ (.CLK(clknet_leaf_1_clk),
    .D(_00604_),
    .Q(\rvsingle.dp.rf.rf[23][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13147_ (.CLK(clknet_leaf_142_clk),
    .D(_00605_),
    .Q(\rvsingle.dp.rf.rf[23][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13148_ (.CLK(clknet_leaf_147_clk),
    .D(_00606_),
    .Q(\rvsingle.dp.rf.rf[23][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13149_ (.CLK(clknet_leaf_143_clk),
    .D(_00607_),
    .Q(\rvsingle.dp.rf.rf[23][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13150_ (.CLK(clknet_leaf_0_clk),
    .D(_00608_),
    .Q(\rvsingle.dp.rf.rf[23][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13151_ (.CLK(clknet_leaf_0_clk),
    .D(_00609_),
    .Q(\rvsingle.dp.rf.rf[23][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13152_ (.CLK(clknet_leaf_118_clk),
    .D(_00610_),
    .Q(\rvsingle.dp.rf.rf[23][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13153_ (.CLK(clknet_leaf_140_clk),
    .D(_00611_),
    .Q(\rvsingle.dp.rf.rf[23][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13154_ (.CLK(clknet_leaf_128_clk),
    .D(_00612_),
    .Q(\rvsingle.dp.rf.rf[23][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13155_ (.CLK(clknet_leaf_118_clk),
    .D(_00613_),
    .Q(\rvsingle.dp.rf.rf[23][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13156_ (.CLK(clknet_leaf_109_clk),
    .D(_00614_),
    .Q(\rvsingle.dp.rf.rf[23][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13157_ (.CLK(clknet_leaf_115_clk),
    .D(_00615_),
    .Q(\rvsingle.dp.rf.rf[23][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13158_ (.CLK(clknet_leaf_113_clk),
    .D(_00616_),
    .Q(\rvsingle.dp.rf.rf[23][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13159_ (.CLK(clknet_leaf_99_clk),
    .D(_00617_),
    .Q(\rvsingle.dp.rf.rf[23][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13160_ (.CLK(clknet_leaf_103_clk),
    .D(_00618_),
    .Q(\rvsingle.dp.rf.rf[23][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13161_ (.CLK(clknet_leaf_95_clk),
    .D(_00619_),
    .Q(\rvsingle.dp.rf.rf[23][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13162_ (.CLK(clknet_leaf_82_clk),
    .D(_00620_),
    .Q(\rvsingle.dp.rf.rf[23][31] ));
 sky130_fd_sc_hd__dfrtp_2 _13163_ (.CLK(clknet_leaf_74_clk),
    .D(_00621_),
    .RESET_B(_00000_),
    .Q(PC[0]));
 sky130_fd_sc_hd__dfrtp_2 _13164_ (.CLK(clknet_leaf_84_clk),
    .D(_00622_),
    .RESET_B(_00001_),
    .Q(PC[1]));
 sky130_fd_sc_hd__dfxtp_2 _13165_ (.CLK(clknet_leaf_90_clk),
    .D(_00623_),
    .Q(\rvsingle.dp.rf.rf[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13166_ (.CLK(clknet_leaf_53_clk),
    .D(_00624_),
    .Q(\rvsingle.dp.rf.rf[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13167_ (.CLK(clknet_leaf_49_clk),
    .D(_00625_),
    .Q(\rvsingle.dp.rf.rf[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13168_ (.CLK(clknet_leaf_71_clk),
    .D(_00626_),
    .Q(\rvsingle.dp.rf.rf[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13169_ (.CLK(clknet_leaf_58_clk),
    .D(_00627_),
    .Q(\rvsingle.dp.rf.rf[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13170_ (.CLK(clknet_leaf_51_clk),
    .D(_00628_),
    .Q(\rvsingle.dp.rf.rf[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13171_ (.CLK(clknet_leaf_48_clk),
    .D(_00629_),
    .Q(\rvsingle.dp.rf.rf[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13172_ (.CLK(clknet_leaf_56_clk),
    .D(_00630_),
    .Q(\rvsingle.dp.rf.rf[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13173_ (.CLK(clknet_leaf_17_clk),
    .D(_00631_),
    .Q(\rvsingle.dp.rf.rf[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13174_ (.CLK(clknet_leaf_62_clk),
    .D(_00632_),
    .Q(\rvsingle.dp.rf.rf[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13175_ (.CLK(clknet_leaf_65_clk),
    .D(_00633_),
    .Q(\rvsingle.dp.rf.rf[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13176_ (.CLK(clknet_leaf_22_clk),
    .D(_00634_),
    .Q(\rvsingle.dp.rf.rf[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13177_ (.CLK(clknet_leaf_16_clk),
    .D(_00635_),
    .Q(\rvsingle.dp.rf.rf[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13178_ (.CLK(clknet_leaf_20_clk),
    .D(_00636_),
    .Q(\rvsingle.dp.rf.rf[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13179_ (.CLK(clknet_leaf_18_clk),
    .D(_00637_),
    .Q(\rvsingle.dp.rf.rf[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13180_ (.CLK(clknet_leaf_14_clk),
    .D(_00638_),
    .Q(\rvsingle.dp.rf.rf[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13181_ (.CLK(clknet_leaf_139_clk),
    .D(_00639_),
    .Q(\rvsingle.dp.rf.rf[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13182_ (.CLK(clknet_leaf_147_clk),
    .D(_00640_),
    .Q(\rvsingle.dp.rf.rf[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13183_ (.CLK(clknet_leaf_144_clk),
    .D(_00641_),
    .Q(\rvsingle.dp.rf.rf[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13184_ (.CLK(clknet_leaf_13_clk),
    .D(_00642_),
    .Q(\rvsingle.dp.rf.rf[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13185_ (.CLK(clknet_leaf_133_clk),
    .D(_00643_),
    .Q(\rvsingle.dp.rf.rf[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13186_ (.CLK(clknet_leaf_138_clk),
    .D(_00644_),
    .Q(\rvsingle.dp.rf.rf[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13187_ (.CLK(clknet_leaf_130_clk),
    .D(_00645_),
    .Q(\rvsingle.dp.rf.rf[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13188_ (.CLK(clknet_leaf_137_clk),
    .D(_00646_),
    .Q(\rvsingle.dp.rf.rf[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13189_ (.CLK(clknet_leaf_125_clk),
    .D(_00647_),
    .Q(\rvsingle.dp.rf.rf[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13190_ (.CLK(clknet_leaf_111_clk),
    .D(_00648_),
    .Q(\rvsingle.dp.rf.rf[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13191_ (.CLK(clknet_leaf_101_clk),
    .D(_00649_),
    .Q(\rvsingle.dp.rf.rf[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13192_ (.CLK(clknet_leaf_121_clk),
    .D(_00650_),
    .Q(\rvsingle.dp.rf.rf[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13193_ (.CLK(clknet_leaf_100_clk),
    .D(_00651_),
    .Q(\rvsingle.dp.rf.rf[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13194_ (.CLK(clknet_leaf_102_clk),
    .D(_00652_),
    .Q(\rvsingle.dp.rf.rf[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13195_ (.CLK(clknet_leaf_92_clk),
    .D(_00653_),
    .Q(\rvsingle.dp.rf.rf[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13196_ (.CLK(clknet_leaf_93_clk),
    .D(_00654_),
    .Q(\rvsingle.dp.rf.rf[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13197_ (.CLK(clknet_leaf_90_clk),
    .D(_00655_),
    .Q(\rvsingle.dp.rf.rf[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13198_ (.CLK(clknet_leaf_53_clk),
    .D(_00656_),
    .Q(\rvsingle.dp.rf.rf[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13199_ (.CLK(clknet_leaf_44_clk),
    .D(_00657_),
    .Q(\rvsingle.dp.rf.rf[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13200_ (.CLK(clknet_leaf_70_clk),
    .D(_00658_),
    .Q(\rvsingle.dp.rf.rf[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13201_ (.CLK(clknet_leaf_55_clk),
    .D(_00659_),
    .Q(\rvsingle.dp.rf.rf[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13202_ (.CLK(clknet_leaf_53_clk),
    .D(_00660_),
    .Q(\rvsingle.dp.rf.rf[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13203_ (.CLK(clknet_leaf_48_clk),
    .D(_00661_),
    .Q(\rvsingle.dp.rf.rf[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13204_ (.CLK(clknet_leaf_55_clk),
    .D(_00662_),
    .Q(\rvsingle.dp.rf.rf[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13205_ (.CLK(clknet_leaf_24_clk),
    .D(_00663_),
    .Q(\rvsingle.dp.rf.rf[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13206_ (.CLK(clknet_leaf_64_clk),
    .D(_00664_),
    .Q(\rvsingle.dp.rf.rf[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13207_ (.CLK(clknet_leaf_64_clk),
    .D(_00665_),
    .Q(\rvsingle.dp.rf.rf[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13208_ (.CLK(clknet_leaf_22_clk),
    .D(_00666_),
    .Q(\rvsingle.dp.rf.rf[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13209_ (.CLK(clknet_leaf_15_clk),
    .D(_00667_),
    .Q(\rvsingle.dp.rf.rf[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13210_ (.CLK(clknet_leaf_21_clk),
    .D(_00668_),
    .Q(\rvsingle.dp.rf.rf[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13211_ (.CLK(clknet_leaf_17_clk),
    .D(_00669_),
    .Q(\rvsingle.dp.rf.rf[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13212_ (.CLK(clknet_leaf_14_clk),
    .D(_00670_),
    .Q(\rvsingle.dp.rf.rf[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13213_ (.CLK(clknet_leaf_139_clk),
    .D(_00671_),
    .Q(\rvsingle.dp.rf.rf[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13214_ (.CLK(clknet_leaf_148_clk),
    .D(_00672_),
    .Q(\rvsingle.dp.rf.rf[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13215_ (.CLK(clknet_leaf_148_clk),
    .D(_00673_),
    .Q(\rvsingle.dp.rf.rf[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13216_ (.CLK(clknet_leaf_132_clk),
    .D(_00674_),
    .Q(\rvsingle.dp.rf.rf[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13217_ (.CLK(clknet_leaf_128_clk),
    .D(_00675_),
    .Q(\rvsingle.dp.rf.rf[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13218_ (.CLK(clknet_leaf_137_clk),
    .D(_00676_),
    .Q(\rvsingle.dp.rf.rf[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13219_ (.CLK(clknet_leaf_125_clk),
    .D(_00677_),
    .Q(\rvsingle.dp.rf.rf[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13220_ (.CLK(clknet_leaf_131_clk),
    .D(_00678_),
    .Q(\rvsingle.dp.rf.rf[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13221_ (.CLK(clknet_leaf_123_clk),
    .D(_00679_),
    .Q(\rvsingle.dp.rf.rf[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13222_ (.CLK(clknet_leaf_91_clk),
    .D(_00680_),
    .Q(\rvsingle.dp.rf.rf[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13223_ (.CLK(clknet_leaf_101_clk),
    .D(_00681_),
    .Q(\rvsingle.dp.rf.rf[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13224_ (.CLK(clknet_leaf_111_clk),
    .D(_00682_),
    .Q(\rvsingle.dp.rf.rf[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13225_ (.CLK(clknet_leaf_127_clk),
    .D(_00683_),
    .Q(\rvsingle.dp.rf.rf[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13226_ (.CLK(clknet_leaf_102_clk),
    .D(_00684_),
    .Q(\rvsingle.dp.rf.rf[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13227_ (.CLK(clknet_leaf_94_clk),
    .D(_00685_),
    .Q(\rvsingle.dp.rf.rf[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13228_ (.CLK(clknet_leaf_93_clk),
    .D(_00686_),
    .Q(\rvsingle.dp.rf.rf[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13229_ (.CLK(clknet_leaf_90_clk),
    .D(_00687_),
    .Q(\rvsingle.dp.rf.rf[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13230_ (.CLK(clknet_leaf_54_clk),
    .D(_00688_),
    .Q(\rvsingle.dp.rf.rf[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13231_ (.CLK(clknet_leaf_45_clk),
    .D(_00689_),
    .Q(\rvsingle.dp.rf.rf[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13232_ (.CLK(clknet_leaf_53_clk),
    .D(_00690_),
    .Q(\rvsingle.dp.rf.rf[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13233_ (.CLK(clknet_leaf_27_clk),
    .D(_00691_),
    .Q(\rvsingle.dp.rf.rf[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13234_ (.CLK(clknet_leaf_55_clk),
    .D(_00692_),
    .Q(\rvsingle.dp.rf.rf[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13235_ (.CLK(clknet_leaf_47_clk),
    .D(_00693_),
    .Q(\rvsingle.dp.rf.rf[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13236_ (.CLK(clknet_leaf_58_clk),
    .D(_00694_),
    .Q(\rvsingle.dp.rf.rf[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13237_ (.CLK(clknet_leaf_10_clk),
    .D(_00695_),
    .Q(\rvsingle.dp.rf.rf[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13238_ (.CLK(clknet_leaf_62_clk),
    .D(_00696_),
    .Q(\rvsingle.dp.rf.rf[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13239_ (.CLK(clknet_leaf_65_clk),
    .D(_00697_),
    .Q(\rvsingle.dp.rf.rf[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13240_ (.CLK(clknet_leaf_24_clk),
    .D(_00698_),
    .Q(\rvsingle.dp.rf.rf[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13241_ (.CLK(clknet_leaf_15_clk),
    .D(_00699_),
    .Q(\rvsingle.dp.rf.rf[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13242_ (.CLK(clknet_leaf_22_clk),
    .D(_00700_),
    .Q(\rvsingle.dp.rf.rf[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13243_ (.CLK(clknet_leaf_10_clk),
    .D(_00701_),
    .Q(\rvsingle.dp.rf.rf[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13244_ (.CLK(clknet_leaf_12_clk),
    .D(_00702_),
    .Q(\rvsingle.dp.rf.rf[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13245_ (.CLK(clknet_leaf_136_clk),
    .D(_00703_),
    .Q(\rvsingle.dp.rf.rf[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13246_ (.CLK(clknet_leaf_147_clk),
    .D(_00704_),
    .Q(\rvsingle.dp.rf.rf[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13247_ (.CLK(clknet_leaf_145_clk),
    .D(_00705_),
    .Q(\rvsingle.dp.rf.rf[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13248_ (.CLK(clknet_leaf_134_clk),
    .D(_00706_),
    .Q(\rvsingle.dp.rf.rf[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13249_ (.CLK(clknet_leaf_128_clk),
    .D(_00707_),
    .Q(\rvsingle.dp.rf.rf[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13250_ (.CLK(clknet_leaf_121_clk),
    .D(_00708_),
    .Q(\rvsingle.dp.rf.rf[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13251_ (.CLK(clknet_leaf_130_clk),
    .D(_00709_),
    .Q(\rvsingle.dp.rf.rf[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13252_ (.CLK(clknet_leaf_19_clk),
    .D(_00710_),
    .Q(\rvsingle.dp.rf.rf[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13253_ (.CLK(clknet_leaf_121_clk),
    .D(_00711_),
    .Q(\rvsingle.dp.rf.rf[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13254_ (.CLK(clknet_leaf_101_clk),
    .D(_00712_),
    .Q(\rvsingle.dp.rf.rf[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13255_ (.CLK(clknet_leaf_110_clk),
    .D(_00713_),
    .Q(\rvsingle.dp.rf.rf[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13256_ (.CLK(clknet_leaf_111_clk),
    .D(_00714_),
    .Q(\rvsingle.dp.rf.rf[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13257_ (.CLK(clknet_leaf_127_clk),
    .D(_00715_),
    .Q(\rvsingle.dp.rf.rf[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13258_ (.CLK(clknet_leaf_102_clk),
    .D(_00716_),
    .Q(\rvsingle.dp.rf.rf[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13259_ (.CLK(clknet_leaf_100_clk),
    .D(_00717_),
    .Q(\rvsingle.dp.rf.rf[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13260_ (.CLK(clknet_leaf_93_clk),
    .D(_00718_),
    .Q(\rvsingle.dp.rf.rf[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13261_ (.CLK(clknet_leaf_90_clk),
    .D(_00719_),
    .Q(\rvsingle.dp.rf.rf[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13262_ (.CLK(clknet_leaf_53_clk),
    .D(_00720_),
    .Q(\rvsingle.dp.rf.rf[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13263_ (.CLK(clknet_leaf_48_clk),
    .D(_00721_),
    .Q(\rvsingle.dp.rf.rf[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13264_ (.CLK(clknet_leaf_67_clk),
    .D(_00722_),
    .Q(\rvsingle.dp.rf.rf[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13265_ (.CLK(clknet_leaf_55_clk),
    .D(_00723_),
    .Q(\rvsingle.dp.rf.rf[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13266_ (.CLK(clknet_leaf_67_clk),
    .D(_00724_),
    .Q(\rvsingle.dp.rf.rf[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13267_ (.CLK(clknet_leaf_67_clk),
    .D(_00725_),
    .Q(\rvsingle.dp.rf.rf[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13268_ (.CLK(clknet_leaf_58_clk),
    .D(_00726_),
    .Q(\rvsingle.dp.rf.rf[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13269_ (.CLK(clknet_leaf_24_clk),
    .D(_00727_),
    .Q(\rvsingle.dp.rf.rf[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13270_ (.CLK(clknet_leaf_62_clk),
    .D(_00728_),
    .Q(\rvsingle.dp.rf.rf[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13271_ (.CLK(clknet_leaf_60_clk),
    .D(_00729_),
    .Q(\rvsingle.dp.rf.rf[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13272_ (.CLK(clknet_leaf_26_clk),
    .D(_00730_),
    .Q(\rvsingle.dp.rf.rf[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13273_ (.CLK(clknet_leaf_15_clk),
    .D(_00731_),
    .Q(\rvsingle.dp.rf.rf[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13274_ (.CLK(clknet_leaf_19_clk),
    .D(_00732_),
    .Q(\rvsingle.dp.rf.rf[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13275_ (.CLK(clknet_leaf_23_clk),
    .D(_00733_),
    .Q(\rvsingle.dp.rf.rf[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13276_ (.CLK(clknet_leaf_129_clk),
    .D(_00734_),
    .Q(\rvsingle.dp.rf.rf[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13277_ (.CLK(clknet_leaf_137_clk),
    .D(_00735_),
    .Q(\rvsingle.dp.rf.rf[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13278_ (.CLK(clknet_leaf_146_clk),
    .D(_00736_),
    .Q(\rvsingle.dp.rf.rf[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13279_ (.CLK(clknet_leaf_135_clk),
    .D(_00737_),
    .Q(\rvsingle.dp.rf.rf[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13280_ (.CLK(clknet_leaf_13_clk),
    .D(_00738_),
    .Q(\rvsingle.dp.rf.rf[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13281_ (.CLK(clknet_leaf_131_clk),
    .D(_00739_),
    .Q(\rvsingle.dp.rf.rf[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13282_ (.CLK(clknet_leaf_119_clk),
    .D(_00740_),
    .Q(\rvsingle.dp.rf.rf[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13283_ (.CLK(clknet_leaf_125_clk),
    .D(_00741_),
    .Q(\rvsingle.dp.rf.rf[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13284_ (.CLK(clknet_leaf_131_clk),
    .D(_00742_),
    .Q(\rvsingle.dp.rf.rf[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13285_ (.CLK(clknet_leaf_124_clk),
    .D(_00743_),
    .Q(\rvsingle.dp.rf.rf[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13286_ (.CLK(clknet_leaf_122_clk),
    .D(_00744_),
    .Q(\rvsingle.dp.rf.rf[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13287_ (.CLK(clknet_leaf_89_clk),
    .D(_00745_),
    .Q(\rvsingle.dp.rf.rf[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13288_ (.CLK(clknet_leaf_121_clk),
    .D(_00746_),
    .Q(\rvsingle.dp.rf.rf[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13289_ (.CLK(clknet_leaf_99_clk),
    .D(_00747_),
    .Q(\rvsingle.dp.rf.rf[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13290_ (.CLK(clknet_leaf_103_clk),
    .D(_00748_),
    .Q(\rvsingle.dp.rf.rf[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13291_ (.CLK(clknet_leaf_100_clk),
    .D(_00749_),
    .Q(\rvsingle.dp.rf.rf[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13292_ (.CLK(clknet_leaf_93_clk),
    .D(_00750_),
    .Q(\rvsingle.dp.rf.rf[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13293_ (.CLK(clknet_leaf_89_clk),
    .D(_00751_),
    .Q(\rvsingle.dp.rf.rf[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13294_ (.CLK(clknet_leaf_53_clk),
    .D(_00752_),
    .Q(\rvsingle.dp.rf.rf[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13295_ (.CLK(clknet_leaf_44_clk),
    .D(_00753_),
    .Q(\rvsingle.dp.rf.rf[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13296_ (.CLK(clknet_leaf_67_clk),
    .D(_00754_),
    .Q(\rvsingle.dp.rf.rf[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13297_ (.CLK(clknet_leaf_59_clk),
    .D(_00755_),
    .Q(\rvsingle.dp.rf.rf[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13298_ (.CLK(clknet_leaf_67_clk),
    .D(_00756_),
    .Q(\rvsingle.dp.rf.rf[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13299_ (.CLK(clknet_leaf_68_clk),
    .D(_00757_),
    .Q(\rvsingle.dp.rf.rf[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13300_ (.CLK(clknet_leaf_58_clk),
    .D(_00758_),
    .Q(\rvsingle.dp.rf.rf[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13301_ (.CLK(clknet_leaf_29_clk),
    .D(_00759_),
    .Q(\rvsingle.dp.rf.rf[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13302_ (.CLK(clknet_leaf_62_clk),
    .D(_00760_),
    .Q(\rvsingle.dp.rf.rf[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13303_ (.CLK(clknet_leaf_60_clk),
    .D(_00761_),
    .Q(\rvsingle.dp.rf.rf[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13304_ (.CLK(clknet_leaf_26_clk),
    .D(_00762_),
    .Q(\rvsingle.dp.rf.rf[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13305_ (.CLK(clknet_leaf_19_clk),
    .D(_00763_),
    .Q(\rvsingle.dp.rf.rf[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13306_ (.CLK(clknet_leaf_19_clk),
    .D(_00764_),
    .Q(\rvsingle.dp.rf.rf[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13307_ (.CLK(clknet_leaf_23_clk),
    .D(_00765_),
    .Q(\rvsingle.dp.rf.rf[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13308_ (.CLK(clknet_leaf_14_clk),
    .D(_00766_),
    .Q(\rvsingle.dp.rf.rf[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13309_ (.CLK(clknet_leaf_137_clk),
    .D(_00767_),
    .Q(\rvsingle.dp.rf.rf[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13310_ (.CLK(clknet_leaf_146_clk),
    .D(_00768_),
    .Q(\rvsingle.dp.rf.rf[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13311_ (.CLK(clknet_leaf_135_clk),
    .D(_00769_),
    .Q(\rvsingle.dp.rf.rf[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13312_ (.CLK(clknet_leaf_133_clk),
    .D(_00770_),
    .Q(\rvsingle.dp.rf.rf[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13313_ (.CLK(clknet_leaf_132_clk),
    .D(_00771_),
    .Q(\rvsingle.dp.rf.rf[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13314_ (.CLK(clknet_leaf_120_clk),
    .D(_00772_),
    .Q(\rvsingle.dp.rf.rf[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13315_ (.CLK(clknet_leaf_126_clk),
    .D(_00773_),
    .Q(\rvsingle.dp.rf.rf[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13316_ (.CLK(clknet_leaf_131_clk),
    .D(_00774_),
    .Q(\rvsingle.dp.rf.rf[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13317_ (.CLK(clknet_leaf_126_clk),
    .D(_00775_),
    .Q(\rvsingle.dp.rf.rf[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13318_ (.CLK(clknet_leaf_124_clk),
    .D(_00776_),
    .Q(\rvsingle.dp.rf.rf[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13319_ (.CLK(clknet_leaf_121_clk),
    .D(_00777_),
    .Q(\rvsingle.dp.rf.rf[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13320_ (.CLK(clknet_leaf_121_clk),
    .D(_00778_),
    .Q(\rvsingle.dp.rf.rf[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13321_ (.CLK(clknet_leaf_99_clk),
    .D(_00779_),
    .Q(\rvsingle.dp.rf.rf[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13322_ (.CLK(clknet_leaf_104_clk),
    .D(_00780_),
    .Q(\rvsingle.dp.rf.rf[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13323_ (.CLK(clknet_leaf_127_clk),
    .D(_00781_),
    .Q(\rvsingle.dp.rf.rf[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13324_ (.CLK(clknet_leaf_93_clk),
    .D(_00782_),
    .Q(\rvsingle.dp.rf.rf[3][31] ));
 sky130_fd_sc_hd__dfrtp_2 _13325_ (.CLK(clknet_4_12_0_clk),
    .D(\rvsingle.dp.PCNext[2] ),
    .RESET_B(_00002_),
    .Q(PC[2]));
 sky130_fd_sc_hd__dfrtp_2 _13326_ (.CLK(clknet_leaf_76_clk),
    .D(\rvsingle.dp.PCNext[3] ),
    .RESET_B(_00003_),
    .Q(PC[3]));
 sky130_fd_sc_hd__dfrtp_2 _13327_ (.CLK(clknet_leaf_76_clk),
    .D(\rvsingle.dp.PCNext[4] ),
    .RESET_B(_00004_),
    .Q(PC[4]));
 sky130_fd_sc_hd__dfrtp_2 _13328_ (.CLK(clknet_leaf_73_clk),
    .D(\rvsingle.dp.PCNext[5] ),
    .RESET_B(_00005_),
    .Q(PC[5]));
 sky130_fd_sc_hd__dfrtp_2 _13329_ (.CLK(clknet_leaf_76_clk),
    .D(\rvsingle.dp.PCNext[6] ),
    .RESET_B(_00006_),
    .Q(PC[6]));
 sky130_fd_sc_hd__dfrtp_2 _13330_ (.CLK(clknet_leaf_73_clk),
    .D(\rvsingle.dp.PCNext[7] ),
    .RESET_B(_00007_),
    .Q(PC[7]));
 sky130_fd_sc_hd__dfrtp_2 _13331_ (.CLK(clknet_leaf_74_clk),
    .D(\rvsingle.dp.PCNext[8] ),
    .RESET_B(_00008_),
    .Q(PC[8]));
 sky130_fd_sc_hd__dfrtp_2 _13332_ (.CLK(clknet_leaf_74_clk),
    .D(\rvsingle.dp.PCNext[9] ),
    .RESET_B(_00009_),
    .Q(PC[9]));
 sky130_fd_sc_hd__dfrtp_2 _13333_ (.CLK(clknet_leaf_76_clk),
    .D(\rvsingle.dp.PCNext[10] ),
    .RESET_B(_00010_),
    .Q(PC[10]));
 sky130_fd_sc_hd__dfrtp_2 _13334_ (.CLK(clknet_leaf_75_clk),
    .D(\rvsingle.dp.PCNext[11] ),
    .RESET_B(_00011_),
    .Q(PC[11]));
 sky130_fd_sc_hd__dfrtp_2 _13335_ (.CLK(clknet_leaf_75_clk),
    .D(\rvsingle.dp.PCNext[12] ),
    .RESET_B(_00012_),
    .Q(PC[12]));
 sky130_fd_sc_hd__dfrtp_2 _13336_ (.CLK(clknet_leaf_75_clk),
    .D(\rvsingle.dp.PCNext[13] ),
    .RESET_B(_00013_),
    .Q(PC[13]));
 sky130_fd_sc_hd__dfrtp_2 _13337_ (.CLK(clknet_leaf_75_clk),
    .D(\rvsingle.dp.PCNext[14] ),
    .RESET_B(_00014_),
    .Q(PC[14]));
 sky130_fd_sc_hd__dfrtp_2 _13338_ (.CLK(clknet_leaf_77_clk),
    .D(\rvsingle.dp.PCNext[15] ),
    .RESET_B(_00015_),
    .Q(PC[15]));
 sky130_fd_sc_hd__dfrtp_2 _13339_ (.CLK(clknet_leaf_77_clk),
    .D(\rvsingle.dp.PCNext[16] ),
    .RESET_B(_00016_),
    .Q(PC[16]));
 sky130_fd_sc_hd__dfrtp_2 _13340_ (.CLK(clknet_leaf_77_clk),
    .D(\rvsingle.dp.PCNext[17] ),
    .RESET_B(_00017_),
    .Q(PC[17]));
 sky130_fd_sc_hd__dfrtp_2 _13341_ (.CLK(clknet_leaf_77_clk),
    .D(\rvsingle.dp.PCNext[18] ),
    .RESET_B(_00018_),
    .Q(PC[18]));
 sky130_fd_sc_hd__dfrtp_2 _13342_ (.CLK(clknet_leaf_84_clk),
    .D(\rvsingle.dp.PCNext[19] ),
    .RESET_B(_00019_),
    .Q(PC[19]));
 sky130_fd_sc_hd__dfrtp_2 _13343_ (.CLK(clknet_leaf_78_clk),
    .D(\rvsingle.dp.PCNext[20] ),
    .RESET_B(_00020_),
    .Q(PC[20]));
 sky130_fd_sc_hd__dfrtp_2 _13344_ (.CLK(clknet_leaf_78_clk),
    .D(\rvsingle.dp.PCNext[21] ),
    .RESET_B(_00021_),
    .Q(PC[21]));
 sky130_fd_sc_hd__dfrtp_2 _13345_ (.CLK(clknet_leaf_79_clk),
    .D(\rvsingle.dp.PCNext[22] ),
    .RESET_B(_00022_),
    .Q(PC[22]));
 sky130_fd_sc_hd__dfrtp_2 _13346_ (.CLK(clknet_leaf_79_clk),
    .D(\rvsingle.dp.PCNext[23] ),
    .RESET_B(_00023_),
    .Q(PC[23]));
 sky130_fd_sc_hd__dfrtp_2 _13347_ (.CLK(clknet_leaf_78_clk),
    .D(\rvsingle.dp.PCNext[24] ),
    .RESET_B(_00024_),
    .Q(PC[24]));
 sky130_fd_sc_hd__dfrtp_2 _13348_ (.CLK(clknet_leaf_78_clk),
    .D(\rvsingle.dp.PCNext[25] ),
    .RESET_B(_00025_),
    .Q(PC[25]));
 sky130_fd_sc_hd__dfrtp_2 _13349_ (.CLK(clknet_leaf_79_clk),
    .D(\rvsingle.dp.PCNext[26] ),
    .RESET_B(_00026_),
    .Q(PC[26]));
 sky130_fd_sc_hd__dfrtp_2 _13350_ (.CLK(clknet_leaf_79_clk),
    .D(\rvsingle.dp.PCNext[27] ),
    .RESET_B(_00027_),
    .Q(PC[27]));
 sky130_fd_sc_hd__dfrtp_2 _13351_ (.CLK(clknet_leaf_79_clk),
    .D(\rvsingle.dp.PCNext[28] ),
    .RESET_B(_00028_),
    .Q(PC[28]));
 sky130_fd_sc_hd__dfrtp_2 _13352_ (.CLK(clknet_leaf_80_clk),
    .D(\rvsingle.dp.PCNext[29] ),
    .RESET_B(_00029_),
    .Q(PC[29]));
 sky130_fd_sc_hd__dfrtp_2 _13353_ (.CLK(clknet_leaf_80_clk),
    .D(\rvsingle.dp.PCNext[30] ),
    .RESET_B(_00030_),
    .Q(PC[30]));
 sky130_fd_sc_hd__dfrtp_2 _13354_ (.CLK(clknet_leaf_80_clk),
    .D(\rvsingle.dp.PCNext[31] ),
    .RESET_B(_00031_),
    .Q(PC[31]));
 sky130_fd_sc_hd__dfxtp_2 _13355_ (.CLK(clknet_leaf_86_clk),
    .D(_00783_),
    .Q(\rvsingle.dp.rf.rf[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13356_ (.CLK(clknet_leaf_67_clk),
    .D(_00784_),
    .Q(\rvsingle.dp.rf.rf[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13357_ (.CLK(clknet_leaf_45_clk),
    .D(_00785_),
    .Q(\rvsingle.dp.rf.rf[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13358_ (.CLK(clknet_leaf_68_clk),
    .D(_00786_),
    .Q(\rvsingle.dp.rf.rf[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13359_ (.CLK(clknet_leaf_66_clk),
    .D(_00787_),
    .Q(\rvsingle.dp.rf.rf[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13360_ (.CLK(clknet_leaf_67_clk),
    .D(_00788_),
    .Q(\rvsingle.dp.rf.rf[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13361_ (.CLK(clknet_leaf_56_clk),
    .D(_00789_),
    .Q(\rvsingle.dp.rf.rf[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13362_ (.CLK(clknet_leaf_56_clk),
    .D(_00790_),
    .Q(\rvsingle.dp.rf.rf[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13363_ (.CLK(clknet_leaf_26_clk),
    .D(_00791_),
    .Q(\rvsingle.dp.rf.rf[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13364_ (.CLK(clknet_4_12_0_clk),
    .D(_00792_),
    .Q(\rvsingle.dp.rf.rf[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13365_ (.CLK(clknet_leaf_64_clk),
    .D(_00793_),
    .Q(\rvsingle.dp.rf.rf[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13366_ (.CLK(clknet_leaf_25_clk),
    .D(_00794_),
    .Q(\rvsingle.dp.rf.rf[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13367_ (.CLK(clknet_leaf_16_clk),
    .D(_00795_),
    .Q(\rvsingle.dp.rf.rf[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13368_ (.CLK(clknet_leaf_20_clk),
    .D(_00796_),
    .Q(\rvsingle.dp.rf.rf[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13369_ (.CLK(clknet_leaf_16_clk),
    .D(_00797_),
    .Q(\rvsingle.dp.rf.rf[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13370_ (.CLK(clknet_leaf_14_clk),
    .D(_00798_),
    .Q(\rvsingle.dp.rf.rf[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13371_ (.CLK(clknet_leaf_138_clk),
    .D(_00799_),
    .Q(\rvsingle.dp.rf.rf[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13372_ (.CLK(clknet_leaf_148_clk),
    .D(_00800_),
    .Q(\rvsingle.dp.rf.rf[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13373_ (.CLK(clknet_leaf_144_clk),
    .D(_00801_),
    .Q(\rvsingle.dp.rf.rf[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13374_ (.CLK(clknet_leaf_14_clk),
    .D(_00802_),
    .Q(\rvsingle.dp.rf.rf[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13375_ (.CLK(clknet_leaf_133_clk),
    .D(_00803_),
    .Q(\rvsingle.dp.rf.rf[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13376_ (.CLK(clknet_leaf_120_clk),
    .D(_00804_),
    .Q(\rvsingle.dp.rf.rf[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13377_ (.CLK(clknet_leaf_125_clk),
    .D(_00805_),
    .Q(\rvsingle.dp.rf.rf[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13378_ (.CLK(clknet_leaf_130_clk),
    .D(_00806_),
    .Q(\rvsingle.dp.rf.rf[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13379_ (.CLK(clknet_leaf_124_clk),
    .D(_00807_),
    .Q(\rvsingle.dp.rf.rf[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13380_ (.CLK(clknet_leaf_91_clk),
    .D(_00808_),
    .Q(\rvsingle.dp.rf.rf[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13381_ (.CLK(clknet_leaf_123_clk),
    .D(_00809_),
    .Q(\rvsingle.dp.rf.rf[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13382_ (.CLK(clknet_leaf_122_clk),
    .D(_00810_),
    .Q(\rvsingle.dp.rf.rf[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13383_ (.CLK(clknet_leaf_100_clk),
    .D(_00811_),
    .Q(\rvsingle.dp.rf.rf[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13384_ (.CLK(clknet_leaf_122_clk),
    .D(_00812_),
    .Q(\rvsingle.dp.rf.rf[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13385_ (.CLK(clknet_leaf_94_clk),
    .D(_00813_),
    .Q(\rvsingle.dp.rf.rf[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13386_ (.CLK(clknet_leaf_82_clk),
    .D(_00814_),
    .Q(\rvsingle.dp.rf.rf[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 _13387_ (.CLK(clknet_leaf_87_clk),
    .D(_00815_),
    .Q(\rvsingle.dp.rf.rf[30][0] ));
 sky130_fd_sc_hd__dfxtp_2 _13388_ (.CLK(clknet_leaf_51_clk),
    .D(_00816_),
    .Q(\rvsingle.dp.rf.rf[30][1] ));
 sky130_fd_sc_hd__dfxtp_2 _13389_ (.CLK(clknet_leaf_46_clk),
    .D(_00817_),
    .Q(\rvsingle.dp.rf.rf[30][2] ));
 sky130_fd_sc_hd__dfxtp_2 _13390_ (.CLK(clknet_leaf_65_clk),
    .D(_00818_),
    .Q(\rvsingle.dp.rf.rf[30][3] ));
 sky130_fd_sc_hd__dfxtp_2 _13391_ (.CLK(clknet_leaf_39_clk),
    .D(_00819_),
    .Q(\rvsingle.dp.rf.rf[30][4] ));
 sky130_fd_sc_hd__dfxtp_2 _13392_ (.CLK(clknet_leaf_55_clk),
    .D(_00820_),
    .Q(\rvsingle.dp.rf.rf[30][5] ));
 sky130_fd_sc_hd__dfxtp_2 _13393_ (.CLK(clknet_leaf_48_clk),
    .D(_00821_),
    .Q(\rvsingle.dp.rf.rf[30][6] ));
 sky130_fd_sc_hd__dfxtp_2 _13394_ (.CLK(clknet_leaf_40_clk),
    .D(_00822_),
    .Q(\rvsingle.dp.rf.rf[30][7] ));
 sky130_fd_sc_hd__dfxtp_2 _13395_ (.CLK(clknet_4_8_0_clk),
    .D(_00823_),
    .Q(\rvsingle.dp.rf.rf[30][8] ));
 sky130_fd_sc_hd__dfxtp_2 _13396_ (.CLK(clknet_leaf_21_clk),
    .D(_00824_),
    .Q(\rvsingle.dp.rf.rf[30][9] ));
 sky130_fd_sc_hd__dfxtp_2 _13397_ (.CLK(clknet_leaf_37_clk),
    .D(_00825_),
    .Q(\rvsingle.dp.rf.rf[30][10] ));
 sky130_fd_sc_hd__dfxtp_2 _13398_ (.CLK(clknet_leaf_31_clk),
    .D(_00826_),
    .Q(\rvsingle.dp.rf.rf[30][11] ));
 sky130_fd_sc_hd__dfxtp_2 _13399_ (.CLK(clknet_leaf_6_clk),
    .D(_00827_),
    .Q(\rvsingle.dp.rf.rf[30][12] ));
 sky130_fd_sc_hd__dfxtp_2 _13400_ (.CLK(clknet_leaf_24_clk),
    .D(_00828_),
    .Q(\rvsingle.dp.rf.rf[30][13] ));
 sky130_fd_sc_hd__dfxtp_2 _13401_ (.CLK(clknet_leaf_32_clk),
    .D(_00829_),
    .Q(\rvsingle.dp.rf.rf[30][14] ));
 sky130_fd_sc_hd__dfxtp_2 _13402_ (.CLK(clknet_leaf_5_clk),
    .D(_00830_),
    .Q(\rvsingle.dp.rf.rf[30][15] ));
 sky130_fd_sc_hd__dfxtp_2 _13403_ (.CLK(clknet_leaf_142_clk),
    .D(_00831_),
    .Q(\rvsingle.dp.rf.rf[30][16] ));
 sky130_fd_sc_hd__dfxtp_2 _13404_ (.CLK(clknet_leaf_147_clk),
    .D(_00832_),
    .Q(\rvsingle.dp.rf.rf[30][17] ));
 sky130_fd_sc_hd__dfxtp_2 _13405_ (.CLK(clknet_leaf_143_clk),
    .D(_00833_),
    .Q(\rvsingle.dp.rf.rf[30][18] ));
 sky130_fd_sc_hd__dfxtp_2 _13406_ (.CLK(clknet_leaf_0_clk),
    .D(_00834_),
    .Q(\rvsingle.dp.rf.rf[30][19] ));
 sky130_fd_sc_hd__dfxtp_2 _13407_ (.CLK(clknet_leaf_1_clk),
    .D(_00835_),
    .Q(\rvsingle.dp.rf.rf[30][20] ));
 sky130_fd_sc_hd__dfxtp_2 _13408_ (.CLK(clknet_leaf_119_clk),
    .D(_00836_),
    .Q(\rvsingle.dp.rf.rf[30][21] ));
 sky130_fd_sc_hd__dfxtp_2 _13409_ (.CLK(clknet_leaf_139_clk),
    .D(_00837_),
    .Q(\rvsingle.dp.rf.rf[30][22] ));
 sky130_fd_sc_hd__dfxtp_2 _13410_ (.CLK(clknet_leaf_130_clk),
    .D(_00838_),
    .Q(\rvsingle.dp.rf.rf[30][23] ));
 sky130_fd_sc_hd__dfxtp_2 _13411_ (.CLK(clknet_leaf_121_clk),
    .D(_00839_),
    .Q(\rvsingle.dp.rf.rf[30][24] ));
 sky130_fd_sc_hd__dfxtp_2 _13412_ (.CLK(clknet_leaf_109_clk),
    .D(_00840_),
    .Q(\rvsingle.dp.rf.rf[30][25] ));
 sky130_fd_sc_hd__dfxtp_2 _13413_ (.CLK(clknet_leaf_112_clk),
    .D(_00841_),
    .Q(\rvsingle.dp.rf.rf[30][26] ));
 sky130_fd_sc_hd__dfxtp_2 _13414_ (.CLK(clknet_leaf_113_clk),
    .D(_00842_),
    .Q(\rvsingle.dp.rf.rf[30][27] ));
 sky130_fd_sc_hd__dfxtp_2 _13415_ (.CLK(clknet_leaf_101_clk),
    .D(_00843_),
    .Q(\rvsingle.dp.rf.rf[30][28] ));
 sky130_fd_sc_hd__dfxtp_2 _13416_ (.CLK(clknet_leaf_106_clk),
    .D(_00844_),
    .Q(\rvsingle.dp.rf.rf[30][29] ));
 sky130_fd_sc_hd__dfxtp_2 _13417_ (.CLK(clknet_leaf_94_clk),
    .D(_00845_),
    .Q(\rvsingle.dp.rf.rf[30][30] ));
 sky130_fd_sc_hd__dfxtp_2 _13418_ (.CLK(clknet_leaf_81_clk),
    .D(_00846_),
    .Q(\rvsingle.dp.rf.rf[30][31] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rvsingle.dp.rf.rf[9][0] ),
    .X(net1));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\rvsingle.dp.rf.rf[25][5] ),
    .X(net2));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\rvsingle.dp.rf.rf[1][9] ),
    .X(net3));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\rvsingle.dp.rf.rf[1][0] ),
    .X(net4));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\rvsingle.dp.rf.rf[25][3] ),
    .X(net5));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\rvsingle.dp.rf.rf[25][20] ),
    .X(net6));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\rvsingle.dp.rf.rf[27][0] ),
    .X(net7));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\rvsingle.dp.rf.rf[24][9] ),
    .X(net8));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\rvsingle.dp.rf.rf[20][0] ),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\rvsingle.dp.rf.rf[25][17] ),
    .X(net10));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\rvsingle.dp.rf.rf[11][7] ),
    .X(net11));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\rvsingle.dp.rf.rf[1][18] ),
    .X(net12));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\rvsingle.dp.rf.rf[1][5] ),
    .X(net13));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\rvsingle.dp.rf.rf[11][9] ),
    .X(net14));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\rvsingle.dp.rf.rf[0][10] ),
    .X(net15));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\rvsingle.dp.rf.rf[16][20] ),
    .X(net16));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\rvsingle.dp.rf.rf[24][0] ),
    .X(net17));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\rvsingle.dp.rf.rf[19][10] ),
    .X(net18));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\rvsingle.dp.rf.rf[3][7] ),
    .X(net19));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\rvsingle.dp.rf.rf[3][18] ),
    .X(net20));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\rvsingle.dp.rf.rf[3][9] ),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\rvsingle.dp.rf.rf[1][16] ),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\rvsingle.dp.rf.rf[24][24] ),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\rvsingle.dp.rf.rf[28][0] ),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\rvsingle.dp.rf.rf[30][31] ),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\rvsingle.dp.rf.rf[27][20] ),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\rvsingle.dp.rf.rf[9][22] ),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\rvsingle.dp.rf.rf[3][0] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\rvsingle.dp.rf.rf[4][31] ),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\rvsingle.dp.rf.rf[27][5] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\rvsingle.dp.rf.rf[11][20] ),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\rvsingle.dp.rf.rf[7][31] ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\rvsingle.dp.rf.rf[0][7] ),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\rvsingle.dp.rf.rf[22][0] ),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\rvsingle.dp.rf.rf[2][0] ),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\rvsingle.dp.rf.rf[7][4] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\rvsingle.dp.rf.rf[7][3] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\rvsingle.dp.rf.rf[12][31] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\rvsingle.dp.rf.rf[1][17] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\rvsingle.dp.rf.rf[22][31] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\rvsingle.dp.rf.rf[28][31] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\rvsingle.dp.rf.rf[27][3] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\rvsingle.dp.rf.rf[6][31] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\rvsingle.dp.rf.rf[23][31] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\rvsingle.dp.rf.rf[5][3] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\rvsingle.dp.rf.rf[16][31] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\rvsingle.dp.rf.rf[20][31] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\rvsingle.dp.rf.rf[10][31] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\rvsingle.dp.rf.rf[8][31] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\rvsingle.dp.rf.rf[9][10] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\rvsingle.dp.rf.rf[19][31] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\rvsingle.dp.rf.rf[5][10] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\rvsingle.dp.rf.rf[30][0] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\rvsingle.dp.rf.rf[17][6] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\rvsingle.dp.rf.rf[11][31] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\rvsingle.dp.rf.rf[18][31] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\rvsingle.dp.rf.rf[17][31] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\rvsingle.dp.rf.rf[21][31] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\rvsingle.dp.rf.rf[13][31] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\rvsingle.dp.rf.rf[11][6] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\rvsingle.dp.rf.rf[0][31] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\rvsingle.dp.rf.rf[3][31] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\rvsingle.dp.rf.rf[19][6] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\rvsingle.dp.rf.rf[9][31] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\rvsingle.dp.rf.rf[19][20] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\rvsingle.dp.rf.rf[9][25] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\rvsingle.dp.rf.rf[25][31] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\rvsingle.dp.rf.rf[27][31] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\rvsingle.dp.rf.rf[7][15] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\rvsingle.dp.rf.rf[15][31] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\rvsingle.dp.rf.rf[14][31] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\rvsingle.dp.rf.rf[19][7] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\rvsingle.dp.rf.rf[1][31] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\rvsingle.dp.rf.rf[29][0] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\rvsingle.dp.rf.rf[25][6] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\rvsingle.dp.rf.rf[11][22] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\rvsingle.dp.rf.rf[24][31] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\rvsingle.dp.rf.rf[9][7] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\rvsingle.dp.rf.rf[7][0] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\rvsingle.dp.rf.rf[29][31] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\rvsingle.dp.rf.rf[31][31] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\rvsingle.dp.rf.rf[5][15] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\rvsingle.dp.rf.rf[5][14] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\rvsingle.dp.rf.rf[26][31] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\rvsingle.dp.rf.rf[3][10] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\rvsingle.dp.rf.rf[11][3] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\rvsingle.dp.rf.rf[19][12] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\rvsingle.dp.rf.rf[9][5] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\rvsingle.dp.rf.rf[5][7] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\rvsingle.dp.rf.rf[5][31] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\rvsingle.dp.rf.rf[7][9] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\rvsingle.dp.rf.rf[7][7] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\rvsingle.dp.rf.rf[11][10] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\rvsingle.dp.rf.rf[9][19] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\rvsingle.dp.rf.rf[7][14] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\rvsingle.dp.rf.rf[5][22] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\rvsingle.dp.rf.rf[3][14] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\rvsingle.dp.rf.rf[1][14] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\rvsingle.dp.rf.rf[2][31] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\rvsingle.dp.rf.rf[3][5] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\rvsingle.dp.rf.rf[7][11] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\rvsingle.dp.rf.rf[11][24] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\rvsingle.dp.rf.rf[3][17] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\rvsingle.dp.rf.rf[11][15] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\rvsingle.dp.rf.rf[7][19] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\rvsingle.dp.rf.rf[27][6] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\rvsingle.dp.rf.rf[19][9] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\rvsingle.dp.rf.rf[17][0] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\rvsingle.dp.rf.rf[19][0] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\rvsingle.dp.rf.rf[16][0] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\rvsingle.dp.rf.rf[6][0] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\rvsingle.dp.rf.rf[31][0] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\rvsingle.dp.rf.rf[11][4] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\rvsingle.dp.rf.rf[9][13] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\rvsingle.dp.rf.rf[18][0] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\rvsingle.dp.rf.rf[4][0] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\rvsingle.dp.rf.rf[7][6] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\rvsingle.dp.rf.rf[1][3] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\rvsingle.dp.rf.rf[7][22] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\rvsingle.dp.rf.rf[23][0] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\rvsingle.dp.rf.rf[17][3] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\rvsingle.dp.rf.rf[17][12] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\rvsingle.dp.rf.rf[16][9] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\rvsingle.dp.rf.rf[14][0] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\rvsingle.dp.rf.rf[11][5] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\rvsingle.dp.rf.rf[19][14] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\rvsingle.dp.rf.rf[21][0] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\rvsingle.dp.rf.rf[5][13] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\rvsingle.dp.rf.rf[5][6] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\rvsingle.dp.rf.rf[25][21] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\rvsingle.dp.rf.rf[19][13] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\rvsingle.dp.rf.rf[1][15] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\rvsingle.dp.rf.rf[19][19] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\rvsingle.dp.rf.rf[5][26] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\rvsingle.dp.rf.rf[17][7] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\rvsingle.dp.rf.rf[12][0] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\rvsingle.dp.rf.rf[17][19] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\rvsingle.dp.rf.rf[3][3] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\rvsingle.dp.rf.rf[9][14] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\rvsingle.dp.rf.rf[19][4] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\rvsingle.dp.rf.rf[3][26] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\rvsingle.dp.rf.rf[15][0] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\rvsingle.dp.rf.rf[11][12] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\rvsingle.dp.rf.rf[27][17] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\rvsingle.dp.rf.rf[1][21] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\rvsingle.dp.rf.rf[25][19] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\rvsingle.dp.rf.rf[0][0] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\rvsingle.dp.rf.rf[26][0] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\rvsingle.dp.rf.rf[8][0] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\rvsingle.dp.rf.rf[9][3] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\rvsingle.dp.rf.rf[3][15] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\rvsingle.dp.rf.rf[8][9] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\rvsingle.dp.rf.rf[7][16] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\rvsingle.dp.rf.rf[27][21] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\rvsingle.dp.rf.rf[9][18] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\rvsingle.dp.rf.rf[27][19] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\rvsingle.dp.rf.rf[11][13] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\rvsingle.dp.rf.rf[17][14] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\rvsingle.dp.rf.rf[17][5] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\rvsingle.dp.rf.rf[11][11] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\rvsingle.dp.rf.rf[8][20] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\rvsingle.dp.rf.rf[17][22] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\rvsingle.dp.rf.rf[11][17] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\rvsingle.dp.rf.rf[5][0] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\rvsingle.dp.rf.rf[7][13] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\rvsingle.dp.rf.rf[24][12] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\rvsingle.dp.rf.rf[17][10] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\rvsingle.dp.rf.rf[8][12] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\rvsingle.dp.rf.rf[1][19] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\rvsingle.dp.rf.rf[5][12] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\rvsingle.dp.rf.rf[5][21] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\rvsingle.dp.rf.rf[11][14] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\rvsingle.dp.rf.rf[19][24] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\rvsingle.dp.rf.rf[3][19] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\rvsingle.dp.rf.rf[11][19] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\rvsingle.dp.rf.rf[3][16] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\rvsingle.dp.rf.rf[3][21] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\rvsingle.dp.rf.rf[13][0] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\rvsingle.dp.rf.rf[17][26] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\rvsingle.dp.rf.rf[0][26] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\rvsingle.dp.rf.rf[5][4] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\rvsingle.dp.rf.rf[4][20] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\rvsingle.dp.rf.rf[17][15] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\rvsingle.dp.rf.rf[1][12] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\rvsingle.dp.rf.rf[11][25] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\rvsingle.dp.rf.rf[9][21] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\rvsingle.dp.rf.rf[10][0] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\rvsingle.dp.rf.rf[17][18] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\rvsingle.dp.rf.rf[19][11] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\rvsingle.dp.rf.rf[7][25] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\rvsingle.dp.rf.rf[17][25] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\rvsingle.dp.rf.rf[3][20] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\rvsingle.dp.rf.rf[1][4] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\rvsingle.dp.rf.rf[3][12] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\rvsingle.dp.rf.rf[1][13] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\rvsingle.dp.rf.rf[19][5] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\rvsingle.dp.rf.rf[16][24] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\rvsingle.dp.rf.rf[17][4] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\rvsingle.dp.rf.rf[19][17] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\rvsingle.dp.rf.rf[19][22] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\rvsingle.dp.rf.rf[3][13] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\rvsingle.dp.rf.rf[19][15] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\rvsingle.dp.rf.rf[3][4] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\rvsingle.dp.rf.rf[19][3] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\rvsingle.dp.rf.rf[1][20] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\rvsingle.dp.rf.rf[1][22] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\rvsingle.dp.rf.rf[3][22] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\rvsingle.dp.rf.rf[17][21] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\rvsingle.dp.rf.rf[7][17] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\rvsingle.dp.rf.rf[1][6] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\rvsingle.dp.rf.rf[3][6] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\rvsingle.dp.rf.rf[9][27] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\rvsingle.dp.rf.rf[19][25] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\rvsingle.dp.rf.rf[9][26] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\rvsingle.dp.rf.rf[5][27] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\rvsingle.dp.rf.rf[24][28] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\rvsingle.dp.rf.rf[19][16] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\rvsingle.dp.rf.rf[8][11] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\rvsingle.dp.rf.rf[0][29] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\rvsingle.dp.rf.rf[16][22] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\rvsingle.dp.rf.rf[30][28] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\rvsingle.dp.rf.rf[12][29] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\rvsingle.dp.rf.rf[2][26] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\rvsingle.dp.rf.rf[3][11] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\rvsingle.dp.rf.rf[4][27] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\rvsingle.dp.rf.rf[30][23] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\rvsingle.dp.rf.rf[2][15] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\rvsingle.dp.rf.rf[2][28] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\rvsingle.dp.rf.rf[26][24] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\rvsingle.dp.rf.rf[6][22] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\rvsingle.dp.rf.rf[5][11] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\rvsingle.dp.rf.rf[5][16] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\rvsingle.dp.rf.rf[2][30] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\rvsingle.dp.rf.rf[25][22] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\rvsingle.dp.rf.rf[23][28] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\rvsingle.dp.rf.rf[25][28] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\rvsingle.dp.rf.rf[24][16] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\rvsingle.dp.rf.rf[1][23] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\rvsingle.dp.rf.rf[4][29] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\rvsingle.dp.rf.rf[6][27] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\rvsingle.dp.rf.rf[4][19] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\rvsingle.dp.rf.rf[8][23] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\rvsingle.dp.rf.rf[4][30] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\rvsingle.dp.rf.rf[1][24] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\rvsingle.dp.rf.rf[25][23] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\rvsingle.dp.rf.rf[23][14] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\rvsingle.dp.rf.rf[8][30] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\rvsingle.dp.rf.rf[11][0] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\rvsingle.dp.rf.rf[6][24] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\rvsingle.dp.rf.rf[19][23] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\rvsingle.dp.rf.rf[7][12] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\rvsingle.dp.rf.rf[4][28] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\rvsingle.dp.rf.rf[12][2] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\rvsingle.dp.rf.rf[9][24] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\rvsingle.dp.rf.rf[11][29] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\rvsingle.dp.rf.rf[23][23] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\rvsingle.dp.rf.rf[19][28] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\rvsingle.dp.rf.rf[30][30] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\rvsingle.dp.rf.rf[10][24] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\rvsingle.dp.rf.rf[6][25] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\rvsingle.dp.rf.rf[30][29] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\rvsingle.dp.rf.rf[4][26] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\rvsingle.dp.rf.rf[12][30] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\rvsingle.dp.rf.rf[5][28] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\rvsingle.dp.rf.rf[0][17] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\rvsingle.dp.rf.rf[23][30] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\rvsingle.dp.rf.rf[0][30] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\rvsingle.dp.rf.rf[30][26] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\rvsingle.dp.rf.rf[23][9] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\rvsingle.dp.rf.rf[23][8] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\rvsingle.dp.rf.rf[18][23] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\rvsingle.dp.rf.rf[27][30] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\rvsingle.dp.rf.rf[28][20] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\rvsingle.dp.rf.rf[27][24] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\rvsingle.dp.rf.rf[4][4] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\rvsingle.dp.rf.rf[5][29] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\rvsingle.dp.rf.rf[7][28] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\rvsingle.dp.rf.rf[4][21] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\rvsingle.dp.rf.rf[28][21] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\rvsingle.dp.rf.rf[1][1] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\rvsingle.dp.rf.rf[10][28] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\rvsingle.dp.rf.rf[12][17] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\rvsingle.dp.rf.rf[26][9] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\rvsingle.dp.rf.rf[30][11] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\rvsingle.dp.rf.rf[19][29] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\rvsingle.dp.rf.rf[28][28] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\rvsingle.dp.rf.rf[10][29] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\rvsingle.dp.rf.rf[8][29] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\rvsingle.dp.rf.rf[27][28] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\rvsingle.dp.rf.rf[17][17] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\rvsingle.dp.rf.rf[29][28] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\rvsingle.dp.rf.rf[6][28] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\rvsingle.dp.rf.rf[4][25] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\rvsingle.dp.rf.rf[9][28] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\rvsingle.dp.rf.rf[14][30] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\rvsingle.dp.rf.rf[1][26] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\rvsingle.dp.rf.rf[26][28] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\rvsingle.dp.rf.rf[23][1] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\rvsingle.dp.rf.rf[11][27] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\rvsingle.dp.rf.rf[1][30] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\rvsingle.dp.rf.rf[28][30] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\rvsingle.dp.rf.rf[29][30] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\rvsingle.dp.rf.rf[5][24] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\rvsingle.dp.rf.rf[2][22] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\rvsingle.dp.rf.rf[30][27] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\rvsingle.dp.rf.rf[28][29] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\rvsingle.dp.rf.rf[3][23] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\rvsingle.dp.rf.rf[25][24] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\rvsingle.dp.rf.rf[12][28] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\rvsingle.dp.rf.rf[7][21] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\rvsingle.dp.rf.rf[17][30] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\rvsingle.dp.rf.rf[9][9] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\rvsingle.dp.rf.rf[3][30] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\rvsingle.dp.rf.rf[4][8] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\rvsingle.dp.rf.rf[26][10] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\rvsingle.dp.rf.rf[5][20] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\rvsingle.dp.rf.rf[23][10] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\rvsingle.dp.rf.rf[21][7] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\rvsingle.dp.rf.rf[1][25] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\rvsingle.dp.rf.rf[26][23] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\rvsingle.dp.rf.rf[4][17] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\rvsingle.dp.rf.rf[27][23] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\rvsingle.dp.rf.rf[24][30] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\rvsingle.dp.rf.rf[3][28] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\rvsingle.dp.rf.rf[21][9] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\rvsingle.dp.rf.rf[21][30] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\rvsingle.dp.rf.rf[4][18] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\rvsingle.dp.rf.rf[29][29] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\rvsingle.dp.rf.rf[6][10] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\rvsingle.dp.rf.rf[22][28] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\rvsingle.dp.rf.rf[0][28] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\rvsingle.dp.rf.rf[19][8] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\rvsingle.dp.rf.rf[23][16] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\rvsingle.dp.rf.rf[9][30] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\rvsingle.dp.rf.rf[16][25] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\rvsingle.dp.rf.rf[6][11] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\rvsingle.dp.rf.rf[26][30] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\rvsingle.dp.rf.rf[12][15] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\rvsingle.dp.rf.rf[2][11] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\rvsingle.dp.rf.rf[18][28] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\rvsingle.dp.rf.rf[24][29] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\rvsingle.dp.rf.rf[1][11] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\rvsingle.dp.rf.rf[25][16] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\rvsingle.dp.rf.rf[20][28] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\rvsingle.dp.rf.rf[21][16] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\rvsingle.dp.rf.rf[10][16] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\rvsingle.dp.rf.rf[22][21] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\rvsingle.dp.rf.rf[0][24] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\rvsingle.dp.rf.rf[18][17] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\rvsingle.dp.rf.rf[27][1] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\rvsingle.dp.rf.rf[16][28] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\rvsingle.dp.rf.rf[7][24] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\rvsingle.dp.rf.rf[26][11] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\rvsingle.dp.rf.rf[4][22] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\rvsingle.dp.rf.rf[31][7] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\rvsingle.dp.rf.rf[0][8] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\rvsingle.dp.rf.rf[8][17] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\rvsingle.dp.rf.rf[8][28] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\rvsingle.dp.rf.rf[7][29] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\rvsingle.dp.rf.rf[6][16] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\rvsingle.dp.rf.rf[16][30] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\rvsingle.dp.rf.rf[0][27] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\rvsingle.dp.rf.rf[10][12] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\rvsingle.dp.rf.rf[18][29] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\rvsingle.dp.rf.rf[21][25] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\rvsingle.dp.rf.rf[26][21] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\rvsingle.dp.rf.rf[13][12] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\rvsingle.dp.rf.rf[12][14] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\rvsingle.dp.rf.rf[22][17] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\rvsingle.dp.rf.rf[25][1] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\rvsingle.dp.rf.rf[25][30] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\rvsingle.dp.rf.rf[9][15] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\rvsingle.dp.rf.rf[30][17] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\rvsingle.dp.rf.rf[17][8] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\rvsingle.dp.rf.rf[4][24] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\rvsingle.dp.rf.rf[2][29] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\rvsingle.dp.rf.rf[6][29] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\rvsingle.dp.rf.rf[3][24] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\rvsingle.dp.rf.rf[10][27] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\rvsingle.dp.rf.rf[13][30] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\rvsingle.dp.rf.rf[8][15] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\rvsingle.dp.rf.rf[26][27] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\rvsingle.dp.rf.rf[1][7] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\rvsingle.dp.rf.rf[6][21] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\rvsingle.dp.rf.rf[18][30] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\rvsingle.dp.rf.rf[4][16] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\rvsingle.dp.rf.rf[12][16] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\rvsingle.dp.rf.rf[3][25] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\rvsingle.dp.rf.rf[25][7] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\rvsingle.dp.rf.rf[8][6] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\rvsingle.dp.rf.rf[2][27] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\rvsingle.dp.rf.rf[23][5] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\rvsingle.dp.rf.rf[28][2] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\rvsingle.dp.rf.rf[28][27] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\rvsingle.dp.rf.rf[12][27] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\rvsingle.dp.rf.rf[8][4] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\rvsingle.dp.rf.rf[10][9] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\rvsingle.dp.rf.rf[0][22] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\rvsingle.dp.rf.rf[16][7] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\rvsingle.dp.rf.rf[4][14] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\rvsingle.dp.rf.rf[30][24] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\rvsingle.dp.rf.rf[22][30] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\rvsingle.dp.rf.rf[2][16] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\rvsingle.dp.rf.rf[29][9] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\rvsingle.dp.rf.rf[26][26] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\rvsingle.dp.rf.rf[2][7] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\rvsingle.dp.rf.rf[15][30] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\rvsingle.dp.rf.rf[17][28] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\rvsingle.dp.rf.rf[8][24] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\rvsingle.dp.rf.rf[14][6] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\rvsingle.dp.rf.rf[21][24] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\rvsingle.dp.rf.rf[10][18] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\rvsingle.dp.rf.rf[20][24] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\rvsingle.dp.rf.rf[6][18] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\rvsingle.dp.rf.rf[28][14] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\rvsingle.dp.rf.rf[26][4] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\rvsingle.dp.rf.rf[26][15] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\rvsingle.dp.rf.rf[26][18] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\rvsingle.dp.rf.rf[29][8] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\rvsingle.dp.rf.rf[2][24] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\rvsingle.dp.rf.rf[28][26] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\rvsingle.dp.rf.rf[10][21] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\rvsingle.dp.rf.rf[21][12] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\rvsingle.dp.rf.rf[20][23] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\rvsingle.dp.rf.rf[26][25] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\rvsingle.dp.rf.rf[31][30] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\rvsingle.dp.rf.rf[14][28] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\rvsingle.dp.rf.rf[0][16] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\rvsingle.dp.rf.rf[16][29] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\rvsingle.dp.rf.rf[21][28] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\rvsingle.dp.rf.rf[29][10] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\rvsingle.dp.rf.rf[16][11] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\rvsingle.dp.rf.rf[6][8] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\rvsingle.dp.rf.rf[28][11] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\rvsingle.dp.rf.rf[5][17] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\rvsingle.dp.rf.rf[24][21] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\rvsingle.dp.rf.rf[2][20] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\rvsingle.dp.rf.rf[15][12] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\rvsingle.dp.rf.rf[5][19] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\rvsingle.dp.rf.rf[15][29] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\rvsingle.dp.rf.rf[19][27] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\rvsingle.dp.rf.rf[11][28] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\rvsingle.dp.rf.rf[31][29] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\rvsingle.dp.rf.rf[29][7] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\rvsingle.dp.rf.rf[24][4] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\rvsingle.dp.rf.rf[26][29] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\rvsingle.dp.rf.rf[20][30] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\rvsingle.dp.rf.rf[17][9] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\rvsingle.dp.rf.rf[15][28] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\rvsingle.dp.rf.rf[0][11] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\rvsingle.dp.rf.rf[16][27] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\rvsingle.dp.rf.rf[10][30] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\rvsingle.dp.rf.rf[24][27] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\rvsingle.dp.rf.rf[21][3] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\rvsingle.dp.rf.rf[31][10] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\rvsingle.dp.rf.rf[26][22] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\rvsingle.dp.rf.rf[26][14] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\rvsingle.dp.rf.rf[14][25] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\rvsingle.dp.rf.rf[14][29] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\rvsingle.dp.rf.rf[16][23] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\rvsingle.dp.rf.rf[20][29] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\rvsingle.dp.rf.rf[24][26] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\rvsingle.dp.rf.rf[20][22] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\rvsingle.dp.rf.rf[28][22] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\rvsingle.dp.rf.rf[13][28] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\rvsingle.dp.rf.rf[8][26] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\rvsingle.dp.rf.rf[12][9] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\rvsingle.dp.rf.rf[14][11] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\rvsingle.dp.rf.rf[26][8] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\rvsingle.dp.rf.rf[8][19] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\rvsingle.dp.rf.rf[17][1] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\rvsingle.dp.rf.rf[0][19] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\rvsingle.dp.rf.rf[14][2] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\rvsingle.dp.rf.rf[5][30] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\rvsingle.dp.rf.rf[30][25] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\rvsingle.dp.rf.rf[8][18] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\rvsingle.dp.rf.rf[23][25] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\rvsingle.dp.rf.rf[9][17] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\rvsingle.dp.rf.rf[22][9] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\rvsingle.dp.rf.rf[25][15] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\rvsingle.dp.rf.rf[30][5] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\rvsingle.dp.rf.rf[0][25] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\rvsingle.dp.rf.rf[19][2] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\rvsingle.dp.rf.rf[13][9] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\rvsingle.dp.rf.rf[20][17] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\rvsingle.dp.rf.rf[11][23] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\rvsingle.dp.rf.rf[6][7] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\rvsingle.dp.rf.rf[13][13] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\rvsingle.dp.rf.rf[1][10] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\rvsingle.dp.rf.rf[30][16] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\rvsingle.dp.rf.rf[18][7] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\rvsingle.dp.rf.rf[6][14] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\rvsingle.dp.rf.rf[10][13] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\rvsingle.dp.rf.rf[5][18] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\rvsingle.dp.rf.rf[14][9] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\rvsingle.dp.rf.rf[25][25] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\rvsingle.dp.rf.rf[7][27] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\rvsingle.dp.rf.rf[23][13] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\rvsingle.dp.rf.rf[21][1] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\rvsingle.dp.rf.rf[21][15] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\rvsingle.dp.rf.rf[15][9] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\rvsingle.dp.rf.rf[31][26] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\rvsingle.dp.rf.rf[13][29] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\rvsingle.dp.rf.rf[28][13] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\rvsingle.dp.rf.rf[23][20] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\rvsingle.dp.rf.rf[30][12] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\rvsingle.dp.rf.rf[22][19] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\rvsingle.dp.rf.rf[15][26] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\rvsingle.dp.rf.rf[13][6] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\rvsingle.dp.rf.rf[18][25] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\rvsingle.dp.rf.rf[3][8] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\rvsingle.dp.rf.rf[14][26] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\rvsingle.dp.rf.rf[0][12] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\rvsingle.dp.rf.rf[22][24] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\rvsingle.dp.rf.rf[28][23] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\rvsingle.dp.rf.rf[10][10] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\rvsingle.dp.rf.rf[20][27] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\rvsingle.dp.rf.rf[19][30] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\rvsingle.dp.rf.rf[2][12] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\rvsingle.dp.rf.rf[6][19] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\rvsingle.dp.rf.rf[21][18] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\rvsingle.dp.rf.rf[16][16] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\rvsingle.dp.rf.rf[25][14] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\rvsingle.dp.rf.rf[2][18] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\rvsingle.dp.rf.rf[30][10] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\rvsingle.dp.rf.rf[6][12] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\rvsingle.dp.rf.rf[8][22] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\rvsingle.dp.rf.rf[24][23] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\rvsingle.dp.rf.rf[18][4] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\rvsingle.dp.rf.rf[8][14] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\rvsingle.dp.rf.rf[0][14] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\rvsingle.dp.rf.rf[0][15] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\rvsingle.dp.rf.rf[16][10] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\rvsingle.dp.rf.rf[29][12] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\rvsingle.dp.rf.rf[9][29] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\rvsingle.dp.rf.rf[23][19] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\rvsingle.dp.rf.rf[8][16] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\rvsingle.dp.rf.rf[2][9] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\rvsingle.dp.rf.rf[24][18] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\rvsingle.dp.rf.rf[0][1] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\rvsingle.dp.rf.rf[11][18] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\rvsingle.dp.rf.rf[6][4] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\rvsingle.dp.rf.rf[6][17] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\rvsingle.dp.rf.rf[15][17] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\rvsingle.dp.rf.rf[26][5] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\rvsingle.dp.rf.rf[22][26] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\rvsingle.dp.rf.rf[7][20] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\rvsingle.dp.rf.rf[21][20] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\rvsingle.dp.rf.rf[4][7] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\rvsingle.dp.rf.rf[10][26] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\rvsingle.dp.rf.rf[0][9] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\rvsingle.dp.rf.rf[10][15] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\rvsingle.dp.rf.rf[6][30] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\rvsingle.dp.rf.rf[0][13] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\rvsingle.dp.rf.rf[18][8] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\rvsingle.dp.rf.rf[12][26] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\rvsingle.dp.rf.rf[18][10] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\rvsingle.dp.rf.rf[22][18] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\rvsingle.dp.rf.rf[13][19] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\rvsingle.dp.rf.rf[4][10] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\rvsingle.dp.rf.rf[6][15] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\rvsingle.dp.rf.rf[23][17] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\rvsingle.dp.rf.rf[19][1] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\rvsingle.dp.rf.rf[11][30] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\rvsingle.dp.rf.rf[27][16] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\rvsingle.dp.rf.rf[12][11] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\rvsingle.dp.rf.rf[22][23] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\rvsingle.dp.rf.rf[23][24] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\rvsingle.dp.rf.rf[12][21] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\rvsingle.dp.rf.rf[2][10] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\rvsingle.dp.rf.rf[20][21] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\rvsingle.dp.rf.rf[16][2] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\rvsingle.dp.rf.rf[26][17] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\rvsingle.dp.rf.rf[30][22] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\rvsingle.dp.rf.rf[22][7] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\rvsingle.dp.rf.rf[4][11] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\rvsingle.dp.rf.rf[18][9] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\rvsingle.dp.rf.rf[8][1] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\rvsingle.dp.rf.rf[6][26] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\rvsingle.dp.rf.rf[27][25] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\rvsingle.dp.rf.rf[25][0] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\rvsingle.dp.rf.rf[2][23] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\rvsingle.dp.rf.rf[20][9] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\rvsingle.dp.rf.rf[10][23] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\rvsingle.dp.rf.rf[8][5] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\rvsingle.dp.rf.rf[25][4] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\rvsingle.dp.rf.rf[10][22] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\rvsingle.dp.rf.rf[7][10] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\rvsingle.dp.rf.rf[20][25] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\rvsingle.dp.rf.rf[14][4] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\rvsingle.dp.rf.rf[20][26] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\rvsingle.dp.rf.rf[9][12] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\rvsingle.dp.rf.rf[30][13] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\rvsingle.dp.rf.rf[18][27] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\rvsingle.dp.rf.rf[17][11] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\rvsingle.dp.rf.rf[5][23] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\rvsingle.dp.rf.rf[26][16] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\rvsingle.dp.rf.rf[10][4] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\rvsingle.dp.rf.rf[30][9] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\rvsingle.dp.rf.rf[28][9] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\rvsingle.dp.rf.rf[26][12] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\rvsingle.dp.rf.rf[2][14] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\rvsingle.dp.rf.rf[29][26] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\rvsingle.dp.rf.rf[14][14] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\rvsingle.dp.rf.rf[2][21] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\rvsingle.dp.rf.rf[17][27] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\rvsingle.dp.rf.rf[8][2] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\rvsingle.dp.rf.rf[0][23] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\rvsingle.dp.rf.rf[22][20] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\rvsingle.dp.rf.rf[30][3] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\rvsingle.dp.rf.rf[13][17] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\rvsingle.dp.rf.rf[28][12] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\rvsingle.dp.rf.rf[8][10] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\rvsingle.dp.rf.rf[18][18] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\rvsingle.dp.rf.rf[2][19] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\rvsingle.dp.rf.rf[25][29] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\rvsingle.dp.rf.rf[11][26] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\rvsingle.dp.rf.rf[14][18] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\rvsingle.dp.rf.rf[21][23] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\rvsingle.dp.rf.rf[5][25] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\rvsingle.dp.rf.rf[29][27] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\rvsingle.dp.rf.rf[30][7] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\rvsingle.dp.rf.rf[12][4] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\rvsingle.dp.rf.rf[22][29] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\rvsingle.dp.rf.rf[24][19] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\rvsingle.dp.rf.rf[24][20] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\rvsingle.dp.rf.rf[12][6] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\rvsingle.dp.rf.rf[12][18] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\rvsingle.dp.rf.rf[0][4] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\rvsingle.dp.rf.rf[21][17] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\rvsingle.dp.rf.rf[12][25] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\rvsingle.dp.rf.rf[10][8] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\rvsingle.dp.rf.rf[16][4] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\rvsingle.dp.rf.rf[18][21] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\rvsingle.dp.rf.rf[23][22] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\rvsingle.dp.rf.rf[5][2] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\rvsingle.dp.rf.rf[31][25] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\rvsingle.dp.rf.rf[1][2] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\rvsingle.dp.rf.rf[27][2] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\rvsingle.dp.rf.rf[13][11] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\rvsingle.dp.rf.rf[1][28] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\rvsingle.dp.rf.rf[0][18] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\rvsingle.dp.rf.rf[6][9] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\rvsingle.dp.rf.rf[31][9] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\rvsingle.dp.rf.rf[13][26] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\rvsingle.dp.rf.rf[15][6] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\rvsingle.dp.rf.rf[20][14] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\rvsingle.dp.rf.rf[2][13] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\rvsingle.dp.rf.rf[7][8] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\rvsingle.dp.rf.rf[21][5] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\rvsingle.dp.rf.rf[30][19] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\rvsingle.dp.rf.rf[17][29] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\rvsingle.dp.rf.rf[12][10] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\rvsingle.dp.rf.rf[17][2] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\rvsingle.dp.rf.rf[4][15] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\rvsingle.dp.rf.rf[28][6] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\rvsingle.dp.rf.rf[31][27] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\rvsingle.dp.rf.rf[16][17] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\rvsingle.dp.rf.rf[25][2] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\rvsingle.dp.rf.rf[7][26] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\rvsingle.dp.rf.rf[23][29] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\rvsingle.dp.rf.rf[22][27] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\rvsingle.dp.rf.rf[12][12] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\rvsingle.dp.rf.rf[9][16] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\rvsingle.dp.rf.rf[6][20] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\rvsingle.dp.rf.rf[8][21] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\rvsingle.dp.rf.rf[3][29] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\rvsingle.dp.rf.rf[29][17] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\rvsingle.dp.rf.rf[9][20] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\rvsingle.dp.rf.rf[21][22] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\rvsingle.dp.rf.rf[9][4] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\rvsingle.dp.rf.rf[22][4] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\rvsingle.dp.rf.rf[16][19] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\rvsingle.dp.rf.rf[0][20] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\rvsingle.dp.rf.rf[23][15] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\rvsingle.dp.rf.rf[2][8] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\rvsingle.dp.rf.rf[8][13] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\rvsingle.dp.rf.rf[24][25] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\rvsingle.dp.rf.rf[4][5] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\rvsingle.dp.rf.rf[4][12] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\rvsingle.dp.rf.rf[12][1] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\rvsingle.dp.rf.rf[12][13] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\rvsingle.dp.rf.rf[21][8] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\rvsingle.dp.rf.rf[3][1] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\rvsingle.dp.rf.rf[20][19] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\rvsingle.dp.rf.rf[12][8] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\rvsingle.dp.rf.rf[2][17] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\rvsingle.dp.rf.rf[30][15] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\rvsingle.dp.rf.rf[31][2] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\rvsingle.dp.rf.rf[11][16] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\rvsingle.dp.rf.rf[23][26] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\rvsingle.dp.rf.rf[17][13] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\rvsingle.dp.rf.rf[25][27] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\rvsingle.dp.rf.rf[22][10] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\rvsingle.dp.rf.rf[12][19] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\rvsingle.dp.rf.rf[23][12] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\rvsingle.dp.rf.rf[13][14] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\rvsingle.dp.rf.rf[31][28] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\rvsingle.dp.rf.rf[7][30] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\rvsingle.dp.rf.rf[30][20] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\rvsingle.dp.rf.rf[14][1] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\rvsingle.dp.rf.rf[16][3] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\rvsingle.dp.rf.rf[6][13] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\rvsingle.dp.rf.rf[1][8] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\rvsingle.dp.rf.rf[29][20] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\rvsingle.dp.rf.rf[30][4] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\rvsingle.dp.rf.rf[28][18] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\rvsingle.dp.rf.rf[14][8] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\rvsingle.dp.rf.rf[31][6] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\rvsingle.dp.rf.rf[27][29] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\rvsingle.dp.rf.rf[22][16] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\rvsingle.dp.rf.rf[18][11] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\rvsingle.dp.rf.rf[13][18] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\rvsingle.dp.rf.rf[7][18] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\rvsingle.dp.rf.rf[11][1] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\rvsingle.dp.rf.rf[30][21] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\rvsingle.dp.rf.rf[15][11] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\rvsingle.dp.rf.rf[26][20] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\rvsingle.dp.rf.rf[10][6] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\rvsingle.dp.rf.rf[13][15] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\rvsingle.dp.rf.rf[23][2] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\rvsingle.dp.rf.rf[27][26] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\rvsingle.dp.rf.rf[13][16] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\rvsingle.dp.rf.rf[15][7] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\rvsingle.dp.rf.rf[14][19] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\rvsingle.dp.rf.rf[13][8] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\rvsingle.dp.rf.rf[8][25] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\rvsingle.dp.rf.rf[14][27] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\rvsingle.dp.rf.rf[15][19] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\rvsingle.dp.rf.rf[27][15] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\rvsingle.dp.rf.rf[24][3] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\rvsingle.dp.rf.rf[28][19] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\rvsingle.dp.rf.rf[26][13] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\rvsingle.dp.rf.rf[6][5] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\rvsingle.dp.rf.rf[22][1] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\rvsingle.dp.rf.rf[12][20] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\rvsingle.dp.rf.rf[31][8] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\rvsingle.dp.rf.rf[24][17] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\rvsingle.dp.rf.rf[20][16] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\rvsingle.dp.rf.rf[29][4] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\rvsingle.dp.rf.rf[15][5] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\rvsingle.dp.rf.rf[28][24] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\rvsingle.dp.rf.rf[10][25] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\rvsingle.dp.rf.rf[15][15] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\rvsingle.dp.rf.rf[22][11] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\rvsingle.dp.rf.rf[18][26] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\rvsingle.dp.rf.rf[22][25] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\rvsingle.dp.rf.rf[28][25] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\rvsingle.dp.rf.rf[30][6] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\rvsingle.dp.rf.rf[21][27] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\rvsingle.dp.rf.rf[4][9] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\rvsingle.dp.rf.rf[29][5] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\rvsingle.dp.rf.rf[13][7] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\rvsingle.dp.rf.rf[22][22] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\rvsingle.dp.rf.rf[28][17] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\rvsingle.dp.rf.rf[21][26] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\rvsingle.dp.rf.rf[29][6] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\rvsingle.dp.rf.rf[23][3] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\rvsingle.dp.rf.rf[2][25] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\rvsingle.dp.rf.rf[30][18] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\rvsingle.dp.rf.rf[14][15] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\rvsingle.dp.rf.rf[26][1] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\rvsingle.dp.rf.rf[27][13] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\rvsingle.dp.rf.rf[25][12] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\rvsingle.dp.rf.rf[24][5] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\rvsingle.dp.rf.rf[29][1] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\rvsingle.dp.rf.rf[9][11] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\rvsingle.dp.rf.rf[9][6] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\rvsingle.dp.rf.rf[25][26] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\rvsingle.dp.rf.rf[24][22] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\rvsingle.dp.rf.rf[24][1] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\rvsingle.dp.rf.rf[31][24] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\rvsingle.dp.rf.rf[21][29] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\rvsingle.dp.rf.rf[28][4] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\rvsingle.dp.rf.rf[3][2] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\rvsingle.dp.rf.rf[14][12] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\rvsingle.dp.rf.rf[8][8] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\rvsingle.dp.rf.rf[23][7] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\rvsingle.dp.rf.rf[23][6] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\rvsingle.dp.rf.rf[23][11] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\rvsingle.dp.rf.rf[18][24] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\rvsingle.dp.rf.rf[20][10] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\rvsingle.dp.rf.rf[21][2] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\rvsingle.dp.rf.rf[23][27] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\rvsingle.dp.rf.rf[14][17] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\rvsingle.dp.rf.rf[26][3] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\rvsingle.dp.rf.rf[25][9] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\rvsingle.dp.rf.rf[15][20] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\rvsingle.dp.rf.rf[26][6] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\rvsingle.dp.rf.rf[20][2] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\rvsingle.dp.rf.rf[0][21] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\rvsingle.dp.rf.rf[8][7] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\rvsingle.dp.rf.rf[16][21] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\rvsingle.dp.rf.rf[20][20] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\rvsingle.dp.rf.rf[16][1] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\rvsingle.dp.rf.rf[29][11] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\rvsingle.dp.rf.rf[27][8] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\rvsingle.dp.rf.rf[2][1] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\rvsingle.dp.rf.rf[7][2] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\rvsingle.dp.rf.rf[29][25] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\rvsingle.dp.rf.rf[13][20] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\rvsingle.dp.rf.rf[22][3] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\rvsingle.dp.rf.rf[15][16] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\rvsingle.dp.rf.rf[30][14] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\rvsingle.dp.rf.rf[29][2] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\rvsingle.dp.rf.rf[15][8] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\rvsingle.dp.rf.rf[20][4] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\rvsingle.dp.rf.rf[7][1] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\rvsingle.dp.rf.rf[28][7] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\rvsingle.dp.rf.rf[14][21] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\rvsingle.dp.rf.rf[23][21] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\rvsingle.dp.rf.rf[31][15] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\rvsingle.dp.rf.rf[19][21] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\rvsingle.dp.rf.rf[8][27] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\rvsingle.dp.rf.rf[31][11] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\rvsingle.dp.rf.rf[29][3] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\rvsingle.dp.rf.rf[18][13] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\rvsingle.dp.rf.rf[25][13] ),
    .X(net818));
endmodule
