
.SUBCKT sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA20 y A1 snd2A1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA21 snd2A1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA20 y A1 snd2A1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA21 snd2A1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB20 pnd2B B1 pndA VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC20 y C1 pnd2B VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA20 y A1 snd2A1 VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA21 snd2A1 A2 VGND VNB nfet_01v8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Y C2 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 net62 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net62 C2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_8 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net36 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net36 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net31 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net35 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net31 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Y A net35 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
rI12 VGND LO sky130_fd_pr__res_generic_po
rI11 HI VPWR sky130_fd_pr__res_generic_po
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net118 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net118 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net181 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net181 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net83 net121 net109 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net109 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net102 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net94 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net94 M1 net102 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net121 clkneg net82 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net83 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net82 net83 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net121 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net166 net83 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net83 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net121 clkpos net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net83 net121 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net145 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net145 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net145 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net83 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net121 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net129 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net80 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net129 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net97 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net89 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net89 S1 net97 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net80 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net141 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net141 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net192 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net192 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net156 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net141 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net141 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net128 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net111 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net96 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net88 S1 net96 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net79 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net111 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net140 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net140 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net191 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net191 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net168 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net168 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net155 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net140 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net140 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=1 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=5 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=5 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net121 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net121 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB special_pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB special_pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net112 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net56 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net112 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net56 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net52 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net52 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net112 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net112 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net107 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net107 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net87 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net87 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net53 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net53 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net44 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net96 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net96 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net76 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net76 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net55 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net55 net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 X net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net55 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net55 net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 X net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
MMIN1 Ab X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 net43 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net43 net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 X net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 net43 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net43 net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net56 net48 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net52 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net48 net44 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net44 net52 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net56 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net56 net48 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net48 net44 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net44 net52 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net52 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
MI14 net124 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net124 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net68 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net92 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net92 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net85 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net85 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net68 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Q_N S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net193 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net193 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net148 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net168 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net168 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net161 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net161 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net148 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net141 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net141 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Q_N S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
MI14 net115 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net115 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net59 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net79 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net83 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net83 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net79 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net76 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net76 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net59 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net175 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net175 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net172 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net160 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net148 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net148 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net172 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net128 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj31 sndNCINn3 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND A sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR A sndPCINp3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 sndPCINp3 CIN majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj31 sndPCINp3 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
MMIN2 COUT net195 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net123 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb mid2 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Bb mid1 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb mid2 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb mid1 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 CIbb CIb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 CIb CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Ab2 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 Abb2 Ab2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 Ab1 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb2 B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab1 Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb2 Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab1 B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT net195 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM net123 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb mid1 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb mid2 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb mid1 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb mid2 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 CIbb CIb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 CIb CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 Ab2 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 Abb2 Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 Ab1 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb2 Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab1 B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb2 B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab1 Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMIP3 SUM net144 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bbb Bb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CINb1 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CINbb2 CINb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CINb2 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CINbb2 mid2 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CINb2 mid1 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bbb mid2 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CINb1 mid1 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net144 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CINb1 mid2 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CINb1 CIN VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CINbb2 CINb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CINb2 CIN VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CINbb2 mid1 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CINb2 mid2 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bbb mid1 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bbb Bb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
MMIP3 SUM net146 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bb2 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb1 mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb1 mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CIb1 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CIbb2 CIb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CIb2 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb1 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb2 mid2 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb2 mid1 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb2 mid2 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb1 mid1 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net146 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb1 mid2 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb1 mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb1 mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CIb1 CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CIbb2 CIb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CIb2 CI VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb1 B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb2 mid1 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb2 mid2 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bb2 mid1 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bb2 B VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_bleeder_1 SHORT VGND VNB VPB VPWR
MI2 net29 SHORT net25 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net25 SHORT net24 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VPWR SHORT net29 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net24 SHORT net16 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net16 SHORT VGND VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_2 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_4 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_8 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_16 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_1 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_2 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_8 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_16 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_3 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_4 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_6 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_8 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_12 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0n_1 A SLEEP_B VGND VNB VPB VPWR X
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net36 A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 sndA SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 net36 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
MI8 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net36 sleepb VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 sleepb SLEEP VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 sleepb sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 sleepb SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 sndA A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1n_1 A SLEEP_B VGND VNB VPB VPWR X
MI23 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 VPWR net44 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 net56 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA net56 net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 net56 SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net44 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X net44 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net44 net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA A net36 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 VPWR net36 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net36 SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputisolatch_1 D SLEEP_B VGND VNB VPB VPWR Q
MI677 Q s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 sleepneg sleeppos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI674 net39 s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 s0 sleepneg net49 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net49 D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 sleeppos net38 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net38 net39 VGND VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 sleeppos SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 sleeppos SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 sleepneg sleeppos VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
MI662 net86 net39 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 sleepneg net86 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net39 s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 s0 sleeppos net69 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net69 D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_16 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 A SLEEP KAPWR VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA net58 net66 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net58 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab net66 KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net66 SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 net66 net58 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net58 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Ab net66 VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 A VGND VPB VPWRIN VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 A LOWLVPWR VGND VNB VPB VPWR X
MI2 net72 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 cross1 net72 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Ab A LOWLVPWR LOWLVPWR pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 X net60 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 net60 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 cross1 Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net72 A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 X net60 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 net60 cross1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 A LOWLVPWR VGND VPB VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
XI1 VGND VNB VPB VPWR net59 LO / sky130_fd_sc_hd__conb_1
XI2 LO LO VGND VNB VPB VPWR nd2right / sky130_fd_sc_hd__nand2_2
XI3 LO LO VGND VNB VPB VPWR nd2left / sky130_fd_sc_hd__nand2_2
XI4 nd2right nd2right VGND VNB VPB VPWR nor2right / sky130_fd_sc_hd__nor2_2
XI5 nd2left nd2left VGND VNB VPB VPWR nor2left / sky130_fd_sc_hd__nor2_2
XI6 nor2right VGND VNB VPB VPWR invright / sky130_fd_sc_hd__inv_2
XI7 nor2left VGND VNB VPB VPWR invleft / sky130_fd_sc_hd__inv_2
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_2 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_4 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA20 VPWR A1 snd2A1 VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA21 snd2A1 A2 y VPB pfet_01v8_hvt w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_0 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.7 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__probe_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net29 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net29 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net29 X sky130_fd_pr__res_generic_m5
.ENDS




.SUBCKT sky130_fd_sc_hd__probec_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net33 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net33 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net33 X short
rI120 VGND met5vgnd short
rI119 VPWR met5vpwr short
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net153 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net153 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net128 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net128 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net103 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net103 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net87 net153 net117 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net117 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net110 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net98 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net98 M1 net110 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net153 clkneg net93 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net87 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net93 net87 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net153 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net87 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net87 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net153 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net87 net153 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net87 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net153 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net83 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net83 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net159 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net159 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net138 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net199 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net199 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net98 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net98 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI27 net243 S1 net215 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net230 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net227 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net199 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net215 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net206 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net199 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net227 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net230 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net243 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net195 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net195 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net130 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net130 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net107 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI34 S0 clkpos net219 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net239 S1 net187 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net230 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net199 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net230 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net219 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net239 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net199 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net195 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net187 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net195 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net212 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net196 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net212 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net196 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net104 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net104 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net177 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net160 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net177 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net160 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net196 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net189 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net196 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net189 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net138 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net123 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net123 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net235 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net235 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net203 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net203 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net240 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net240 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net180 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net180 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net103 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net103 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net179 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net179 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net135 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net135 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net227 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net227 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net206 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net190 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB special_nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net190 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net163 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net163 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd2_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_1 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_2 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_4 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_1 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_2 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_4 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS








































































































































































































.subckt top DataAdr[0] DataAdr[10] DataAdr[11] DataAdr[12] DataAdr[13] DataAdr[14]
+ DataAdr[15] DataAdr[16] DataAdr[17] DataAdr[18] DataAdr[19] DataAdr[1] DataAdr[20]
+ DataAdr[21] DataAdr[22] DataAdr[23] DataAdr[24] DataAdr[25] DataAdr[26] DataAdr[27]
+ DataAdr[28] DataAdr[29] DataAdr[2] DataAdr[30] DataAdr[31] DataAdr[3] DataAdr[4]
+ DataAdr[5] DataAdr[6] DataAdr[7] DataAdr[8] DataAdr[9] Instr[0] Instr[10] Instr[11]
+ Instr[12] Instr[13] Instr[14] Instr[15] Instr[16] Instr[17] Instr[18] Instr[19]
+ Instr[1] Instr[20] Instr[21] Instr[22] Instr[23] Instr[24] Instr[25] Instr[26] Instr[27]
+ Instr[28] Instr[29] Instr[2] Instr[30] Instr[31] Instr[3] Instr[4] Instr[5] Instr[6]
+ Instr[7] Instr[8] Instr[9] MemWrite PC[0] PC[10] PC[11] PC[12] PC[13] PC[14] PC[15]
+ PC[16] PC[17] PC[18] PC[19] PC[1] PC[20] PC[21] PC[22] PC[23] PC[24] PC[25] PC[26]
+ PC[27] PC[28] PC[29] PC[2] PC[30] PC[31] PC[3] PC[4] PC[5] PC[6] PC[7] PC[8] PC[9]
+ ReadData[0] ReadData[10] ReadData[11] ReadData[12] ReadData[13] ReadData[14] ReadData[15]
+ ReadData[16] ReadData[17] ReadData[18] ReadData[19] ReadData[1] ReadData[20] ReadData[21]
+ ReadData[22] ReadData[23] ReadData[24] ReadData[25] ReadData[26] ReadData[27] ReadData[28]
+ ReadData[29] ReadData[2] ReadData[30] ReadData[31] ReadData[3] ReadData[4] ReadData[5]
+ ReadData[6] ReadData[7] ReadData[8] ReadData[9] VGND VPWR WriteData[0] WriteData[10]
+ WriteData[11] WriteData[12] WriteData[13] WriteData[14] WriteData[15] WriteData[16]
+ WriteData[17] WriteData[18] WriteData[19] WriteData[1] WriteData[20] WriteData[21]
+ WriteData[22] WriteData[23] WriteData[24] WriteData[25] WriteData[26] WriteData[27]
+ WriteData[28] WriteData[29] WriteData[2] WriteData[30] WriteData[31] WriteData[3]
+ WriteData[4] WriteData[5] WriteData[6] WriteData[7] WriteData[8] WriteData[9] clk
+ reset
X_06883_ _01591_ _01580_ _01803_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__and3_2
X_09671_ Instr[13] _02912_ _04506_ _04507_ PC[13] VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__a311o_1
X_08622_ _01567_ rvsingle.dp.rf.rf\[16\]\[12\] VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08553_ rvsingle.dp.rf.rf\[0\]\[13\] rvsingle.dp.rf.rf\[1\]\[13\] rvsingle.dp.rf.rf\[2\]\[13\]
+ rvsingle.dp.rf.rf\[3\]\[13\] _01241_ _01953_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__mux4_2
XFILLER_0_77_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07504_ _01156_ _02419_ _02424_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__nand3_1
X_08484_ _03402_ _03403_ _03404_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__nand3_2
XFILLER_0_147_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07435_ _01630_ rvsingle.dp.rf.rf\[30\]\[7\] _01259_ _02355_ VGND VGND VPWR VPWR
+ _02356_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_147_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07366_ rvsingle.dp.rf.rf\[5\]\[7\] _01901_ _02285_ _02286_ VGND VGND VPWR VPWR _02287_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_162_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09105_ _01257_ rvsingle.dp.rf.rf\[8\]\[26\] VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06317_ _01190_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__buf_8
X_07297_ rvsingle.dp.rf.rf\[21\]\[16\] _01513_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__or2b_1
XFILLER_0_45_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09036_ _03943_ _03948_ _01147_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06248_ _01169_ Instr[4] _01170_ Instr[31] VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__o31a_4
XFILLER_0_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold340 rvsingle.dp.rf.rf\[18\]\[28\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06179_ Instr[21] VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold351 rvsingle.dp.rf.rf\[16\]\[28\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 rvsingle.dp.rf.rf\[0\]\[27\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold373 rvsingle.dp.rf.rf\[30\]\[17\] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 rvsingle.dp.rf.rf\[6\]\[21\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 rvsingle.dp.rf.rf\[12\]\[27\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
X_09938_ _04760_ rvsingle.dp.rf.rf\[2\]\[4\] _04741_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__mux2_1
X_09869_ _04693_ _04694_ _04696_ _04697_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__a22o_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _05744_ net336 _05913_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12880_ clknet_leaf_52_clk _00338_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _05000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _04801_ net498 _05874_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__mux2_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _05775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_257 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _05840_ net91 _05742_ _05841_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__a22o_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 _02288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10713_ _05260_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _05805_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10644_ _04863_ net514 _05219_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10575_ _05144_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__buf_4
X_13363_ clknet_leaf_26_clk _00791_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12314_ _04781_ net599 _06099_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13294_ clknet_leaf_53_clk _00752_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12245_ _06074_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__buf_8
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12176_ net176 _06049_ _05345_ _04985_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__a22o_1
X_11127_ _05498_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11058_ _05113_ _05114_ _05115_ _05061_ _04759_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__o311a_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10009_ _04819_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07220_ rvsingle.dp.rf.rf\[5\]\[17\] _01865_ _01668_ _02140_ VGND VGND VPWR VPWR
+ _02141_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07151_ _01688_ rvsingle.dp.rf.rf\[7\]\[18\] _01301_ _02071_ VGND VGND VPWR VPWR
+ _02072_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07082_ _01614_ rvsingle.dp.rf.rf\[6\]\[19\] VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07984_ _02902_ _01617_ _02904_ _02491_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__a31o_1
X_09723_ PC[14] PC[15] PC[16] _04522_ PC[17] VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__a41o_1
X_06935_ _01092_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__clkbuf_8
X_09654_ _04500_ _04501_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__nor2_1
X_06866_ _01783_ _01784_ _01632_ _01786_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__o211ai_1
X_08605_ _01780_ rvsingle.dp.rf.rf\[4\]\[12\] VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nor2_1
X_06797_ _01707_ rvsingle.dp.rf.rf\[18\]\[20\] VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__or2_1
X_09585_ Instr[26] PC[6] VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__xor2_1
XFILLER_0_167_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _01711_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08467_ _02543_ _03385_ _03387_ _01217_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_108_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07418_ _01780_ rvsingle.dp.rf.rf\[2\]\[7\] _02337_ _02338_ VGND VGND VPWR VPWR _02339_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08398_ _02030_ rvsingle.dp.rf.rf\[8\]\[9\] _01104_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_162_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07349_ _01695_ rvsingle.dp.rf.rf\[14\]\[7\] VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10360_ _04721_ _04970_ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__and3_2
XFILLER_0_131_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09019_ _03917_ _03923_ _01248_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__o211ai_4
X_10291_ _04965_ _04927_ _04976_ _04727_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__or4b_4
XFILLER_0_130_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12030_ _04773_ net792 _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold170 rvsingle.dp.rf.rf\[5\]\[12\] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 rvsingle.dp.rf.rf\[5\]\[4\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 rvsingle.dp.rf.rf\[3\]\[20\] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ clknet_leaf_110_clk _00390_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ clknet_leaf_1_clk _00321_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _05534_ net392 _05863_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__mux2_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12794_ clknet_leaf_13_clk _00252_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__buf_4
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11676_ _05728_ rvsingle.dp.rf.rf\[10\]\[2\] _05795_ VGND VGND VPWR VPWR _05797_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13415_ clknet_leaf_101_clk _00843_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10627_ _04818_ net711 _05205_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13346_ clknet_leaf_79_clk rvsingle.dp.PCNext\[23\] _00023_ VGND VGND VPWR VPWR PC[23]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10558_ net155 _05155_ _05174_ _05157_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13277_ clknet_leaf_137_clk _00735_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10489_ _04862_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__buf_2
X_12228_ _06069_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12159_ _05004_ _05324_ _06052_ net138 VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06720_ _01593_ _01624_ _01640_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__nand3_2
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06651_ rvsingle.dp.rf.rf\[7\]\[21\] _01562_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__and2b_1
X_09370_ _01375_ _01406_ _04285_ _04247_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__a211o_2
X_06582_ _01502_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__buf_8
XFILLER_0_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08321_ _03238_ _03239_ _03240_ _03241_ _02483_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08252_ rvsingle.dp.rf.rf\[11\]\[10\] _01677_ _02320_ VGND VGND VPWR VPWR _03173_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07203_ _02120_ _02121_ _01503_ _02123_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08183_ _01630_ rvsingle.dp.rf.rf\[10\]\[11\] VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07134_ rvsingle.dp.rf.rf\[15\]\[18\] _01509_ _02054_ VGND VGND VPWR VPWR _02055_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07065_ _01603_ rvsingle.dp.rf.rf\[8\]\[19\] VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07967_ rvsingle.dp.rf.rf\[30\]\[0\] _01642_ _01596_ VGND VGND VPWR VPWR _02888_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09706_ PC[15] _04536_ _04548_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a21o_1
X_06918_ _01838_ _01804_ _01834_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__o21bai_1
X_07898_ _02815_ _02816_ _02818_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__o21ai_2
X_09637_ _04462_ _04464_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__a21oi_1
X_06849_ rvsingle.dp.rf.rf\[3\]\[23\] _01769_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__or2b_1
XFILLER_0_168_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09568_ _04363_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_167_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08519_ _03434_ _02491_ _03439_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09499_ _03111_ VGND VGND VPWR VPWR WriteData[11] sky130_fd_sc_hd__inv_4
XFILLER_0_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11530_ _05718_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11461_ _05679_ _05643_ _05680_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13200_ clknet_leaf_70_clk _00658_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10412_ _05087_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__clkbuf_1
X_11392_ _04916_ _04918_ _04922_ _05058_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__and4b_2
XFILLER_0_61_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13131_ clknet_leaf_87_clk _00589_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10343_ _04870_ net425 _05044_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13062_ clknet_leaf_113_clk _00520_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10274_ _05011_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12013_ _05099_ _05146_ net149 VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12915_ clknet_leaf_34_clk _00373_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12846_ clknet_leaf_71_clk _00304_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12777_ clknet_leaf_95_clk _00235_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _05713_ net379 _05817_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11659_ _05786_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13329_ clknet_leaf_76_clk rvsingle.dp.PCNext\[6\] _00006_ VGND VGND VPWR VPWR PC[6]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08870_ rvsingle.dp.rf.rf\[12\]\[24\] rvsingle.dp.rf.rf\[13\]\[24\] rvsingle.dp.rf.rf\[14\]\[24\]
+ rvsingle.dp.rf.rf\[15\]\[24\] _01656_ _01260_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07821_ _01650_ rvsingle.dp.rf.rf\[18\]\[3\] _01104_ _02741_ VGND VGND VPWR VPWR
+ _02742_ sky130_fd_sc_hd__o211ai_1
X_07752_ rvsingle.dp.rf.rf\[4\]\[3\] rvsingle.dp.rf.rf\[5\]\[3\] rvsingle.dp.rf.rf\[6\]\[3\]
+ rvsingle.dp.rf.rf\[7\]\[3\] _01903_ _01470_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__mux4_1
X_06703_ _01601_ _01609_ _01116_ _01623_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__o211ai_2
X_07683_ _01687_ rvsingle.dp.rf.rf\[19\]\[5\] _01455_ _02603_ VGND VGND VPWR VPWR
+ _02604_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_126_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09422_ _04325_ _04330_ _04135_ _04331_ VGND VGND VPWR VPWR DataAdr[8] sky130_fd_sc_hd__a31o_4
X_06634_ _01549_ _01550_ _01132_ _01554_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09353_ _01185_ _02261_ _03646_ _03649_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06565_ _01485_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08304_ Instr[30] _01481_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09284_ _03939_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__inv_2
X_06496_ _01416_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08235_ _01725_ rvsingle.dp.rf.rf\[12\]\[10\] VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08166_ _03075_ _01146_ _03086_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__nand3_4
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07117_ rvsingle.dp.rf.rf\[23\]\[18\] _01865_ _02037_ VGND VGND VPWR VPWR _02038_
+ sky130_fd_sc_hd__o21ai_1
X_08097_ _03012_ _02491_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__nand3_1
XFILLER_0_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07048_ _01088_ rvsingle.dp.rf.rf\[21\]\[19\] _01968_ VGND VGND VPWR VPWR _01969_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08999_ rvsingle.dp.rf.rf\[16\]\[27\] rvsingle.dp.rf.rf\[17\]\[27\] _01193_ VGND
+ VGND VPWR VPWR _03919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10961_ _05307_ net594 _05401_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__mux2_1
X_12700_ clknet_leaf_146_clk _00158_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10892_ _04917_ _04965_ _04915_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_38_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12631_ clknet_leaf_6_clk _00089_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12562_ clknet_leaf_59_clk _01046_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11513_ _05352_ rvsingle.dp.rf.rf\[12\]\[23\] _05706_ VGND VGND VPWR VPWR _05709_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12493_ clknet_leaf_44_clk _00977_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11444_ _05671_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11375_ _05633_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13114_ clknet_leaf_14_clk _00572_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10326_ _04824_ net573 _05033_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__mux2_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ clknet_leaf_58_clk _00503_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_10257_ _04828_ rvsingle.dp.rf.rf\[27\]\[18\] _05001_ VGND VGND VPWR VPWR _05002_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10188_ _04957_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12829_ clknet_leaf_143_clk _00287_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06350_ _01157_ _01263_ _01272_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06281_ rvsingle.dp.rf.rf\[12\]\[30\] rvsingle.dp.rf.rf\[13\]\[30\] rvsingle.dp.rf.rf\[14\]\[30\]
+ rvsingle.dp.rf.rf\[15\]\[30\] _01196_ _01203_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_150_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_150_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08020_ _02876_ _01691_ _02940_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold703 rvsingle.dp.rf.rf\[6\]\[13\] VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold714 rvsingle.dp.rf.rf\[7\]\[18\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold725 rvsingle.dp.rf.rf\[14\]\[19\] VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold736 rvsingle.dp.rf.rf\[12\]\[20\] VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold747 rvsingle.dp.rf.rf\[22\]\[25\] VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold758 rvsingle.dp.rf.rf\[23\]\[3\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 rvsingle.dp.rf.rf\[25\]\[26\] VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09971_ _04787_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
X_08922_ _03782_ _03833_ _03835_ _01117_ _03842_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_110_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08853_ _03769_ _03771_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07804_ _01753_ rvsingle.dp.rf.rf\[30\]\[3\] _01596_ _02724_ VGND VGND VPWR VPWR
+ _02725_ sky130_fd_sc_hd__o211ai_2
X_08784_ _01445_ _03700_ _01447_ _03704_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_79_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ _02647_ _02650_ _02364_ _02655_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__o211ai_2
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07666_ rvsingle.dp.rf.rf\[8\]\[5\] rvsingle.dp.rf.rf\[9\]\[5\] _01426_ VGND VGND
+ VPWR VPWR _02587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09405_ _04263_ _04222_ _04135_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__o21ai_2
X_06617_ _01383_ rvsingle.dp.rf.rf\[14\]\[21\] VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07597_ rvsingle.dp.rf.rf\[31\]\[4\] _02481_ _02320_ VGND VGND VPWR VPWR _02518_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09336_ _04250_ _04251_ _02184_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_118_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06548_ _01468_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09267_ _04184_ VGND VGND VPWR VPWR DataAdr[29] sky130_fd_sc_hd__inv_6
XFILLER_0_117_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_141_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_141_clk sky130_fd_sc_hd__clkbuf_16
X_06479_ rvsingle.dp.rf.rf\[8\]\[28\] rvsingle.dp.rf.rf\[9\]\[28\] _01257_ VGND VGND
+ VPWR VPWR _01401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08218_ _01447_ _03131_ _03138_ _02315_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_133_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09198_ Instr[12] Instr[14] _01063_ Instr[13] VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__or4b_4
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08149_ _01382_ rvsingle.dp.rf.rf\[20\]\[11\] VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11160_ _05352_ net460 _05511_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__mux2_1
X_10111_ _04711_ _04743_ _04710_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__and3_1
X_11091_ _05352_ rvsingle.dp.rf.rf\[17\]\[23\] _05469_ VGND VGND VPWR VPWR _05479_
+ sky130_fd_sc_hd__mux2_1
X_10042_ _04846_ net605 _04847_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__mux2_1
Xhold30 rvsingle.dp.rf.rf\[27\]\[5\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 rvsingle.dp.rf.rf\[28\]\[31\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 rvsingle.dp.rf.rf\[5\]\[10\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold63 rvsingle.dp.rf.rf\[19\]\[6\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 rvsingle.dp.rf.rf\[29\]\[0\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 rvsingle.dp.rf.rf\[3\]\[10\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 rvsingle.dp.rf.rf\[5\]\[22\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ _05963_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10944_ _05398_ rvsingle.dp.rf.rf\[18\]\[20\] _05387_ VGND VGND VPWR VPWR _05399_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10875_ _04870_ _05183_ _05336_ _05356_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12614_ clknet_leaf_113_clk _00072_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12545_ clknet_leaf_141_clk _01029_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_132_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_132_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_164_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12476_ clknet_leaf_151_clk _00960_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11427_ _05662_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_5 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11358_ _05624_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10309_ _04782_ net283 _05022_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__mux2_1
X_11289_ _05476_ net544 _05580_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ clknet_leaf_124_clk _00486_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07520_ rvsingle.dp.rf.rf\[0\]\[6\] rvsingle.dp.rf.rf\[1\]\[6\] rvsingle.dp.rf.rf\[2\]\[6\]
+ rvsingle.dp.rf.rf\[3\]\[6\] _02440_ _01470_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07451_ _01152_ _02346_ _02371_ _01083_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__nand4_4
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06402_ _01224_ _01292_ _01314_ _01317_ _01323_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_29_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07382_ _01294_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__clkbuf_8
X_09121_ _04037_ _04038_ _01132_ _04040_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06333_ _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_123_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_123_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09052_ rvsingle.dp.rf.rf\[13\]\[27\] _03857_ _01856_ _03971_ VGND VGND VPWR VPWR
+ _03972_ sky130_fd_sc_hd__o211ai_1
X_06264_ Instr[19] VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__buf_12
XFILLER_0_163_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08003_ rvsingle.dp.rf.rf\[29\]\[0\] _01423_ _01307_ _02923_ VGND VGND VPWR VPWR
+ _02924_ sky130_fd_sc_hd__o211ai_1
Xhold500 rvsingle.dp.rf.rf\[21\]\[15\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
X_06195_ _01102_ _01109_ _01114_ _01118_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold511 rvsingle.dp.rf.rf\[3\]\[8\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold522 rvsingle.dp.rf.rf\[16\]\[16\] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold533 rvsingle.dp.rf.rf\[16\]\[10\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold544 rvsingle.dp.rf.rf\[15\]\[17\] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold555 rvsingle.dp.rf.rf\[18\]\[8\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 rvsingle.dp.rf.rf\[12\]\[11\] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 rvsingle.dp.rf.rf\[18\]\[9\] VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold588 rvsingle.dp.rf.rf\[7\]\[10\] VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ _04773_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__clkbuf_4
Xhold599 rvsingle.dp.rf.rf\[30\]\[9\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ _01184_ _01179_ _03802_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__or3_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _04367_ _04709_ _04712_ _04365_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[31\]
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _03740_ _03744_ _03755_ _03572_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__a41oi_2
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08767_ _02478_ rvsingle.dp.rf.rf\[3\]\[15\] _01490_ _03687_ VGND VGND VPWR VPWR
+ _03688_ sky130_fd_sc_hd__o211ai_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _01743_ rvsingle.dp.rf.rf\[24\]\[5\] VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__nor2_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08698_ _01853_ _03613_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07649_ _01246_ _02550_ _02569_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10660_ _05230_ _05191_ _05231_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09319_ _04210_ _04229_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_114_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_114_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10591_ _04917_ _04727_ _04922_ _04915_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_63_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ _06116_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12261_ _05169_ _05847_ _06077_ net83 VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_120_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11212_ _05391_ rvsingle.dp.rf.rf\[29\]\[14\] _05541_ VGND VGND VPWR VPWR _05545_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12192_ _04885_ rvsingle.dp.rf.rf\[3\]\[27\] _06048_ VGND VGND VPWR VPWR _06062_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11143_ _05212_ rvsingle.dp.rf.rf\[16\]\[15\] _05499_ VGND VGND VPWR VPWR _05507_
+ sky130_fd_sc_hd__mux2_1
X_11074_ _05471_ _05472_ _05463_ net122 VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__a2bb2o_1
X_10025_ _04425_ _04831_ _04832_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a21o_4
XFILLER_0_99_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11976_ _04807_ net400 _05949_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10927_ _05389_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10858_ _05173_ _04726_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__and2_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_105_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10789_ _05303_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__clkbuf_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12528_ clknet_leaf_70_clk _01012_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12459_ clknet_leaf_87_clk _00943_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06951_ rvsingle.dp.rf.rf\[31\]\[22\] _01865_ _01655_ VGND VGND VPWR VPWR _01872_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09670_ _04507_ _04515_ PC[13] VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__o21a_1
X_06882_ _01592_ _01774_ _01802_ _01481_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__nand4_2
X_08621_ _03540_ _03541_ _01511_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08552_ _01694_ _03468_ _01221_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_89_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07503_ _01552_ _02420_ _02421_ _02323_ _02423_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__o311ai_1
X_08483_ _01960_ _02102_ _03318_ _03365_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_77_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07434_ rvsingle.dp.rf.rf\[31\]\[7\] _01566_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07365_ _01725_ rvsingle.dp.rf.rf\[4\]\[7\] VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09104_ rvsingle.dp.rf.rf\[12\]\[26\] rvsingle.dp.rf.rf\[13\]\[26\] rvsingle.dp.rf.rf\[14\]\[26\]
+ rvsingle.dp.rf.rf\[15\]\[26\] _01098_ _03840_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__mux4_1
X_06316_ _01224_ _01228_ _01234_ _01189_ _01238_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07296_ _02213_ _02214_ _01132_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09035_ _01133_ _03949_ _03954_ _01117_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06247_ _01071_ _01079_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__nand2_4
Xhold330 rvsingle.dp.rf.rf\[22\]\[28\] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 rvsingle.dp.rf.rf\[24\]\[29\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ rvsingle.dp.rf.rf\[5\]\[30\] _01090_ _01094_ _01101_ VGND VGND VPWR VPWR
+ _01102_ sky130_fd_sc_hd__o211ai_1
Xhold352 rvsingle.dp.rf.rf\[7\]\[24\] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold363 rvsingle.dp.rf.rf\[10\]\[12\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold374 rvsingle.dp.rf.rf\[17\]\[8\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 rvsingle.dp.rf.rf\[18\]\[30\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 rvsingle.dp.rf.rf\[8\]\[4\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
X_09937_ _04759_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__buf_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ PC[28] PC[29] _04618_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__o21ai_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _03738_ _03739_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__nor2_1
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _04632_ _04633_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__nand2_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _04827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ _05876_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__clkbuf_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_225 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _05841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 DataAdr[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _05843_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__clkbuf_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_269 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10712_ _04859_ net619 _05257_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__mux2_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11692_ _05385_ net516 _05795_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10643_ _05222_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13362_ clknet_leaf_56_clk _00790_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10574_ net214 _05152_ _05182_ _05157_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12313_ _06107_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13293_ clknet_leaf_89_clk _00751_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12244_ _06076_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12175_ _05004_ _05343_ _06052_ net151 VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_102_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11126_ _05381_ net399 _05490_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11057_ _05463_ net121 _05156_ _05464_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10008_ _04818_ net403 _04791_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11959_ _05496_ rvsingle.dp.rf.rf\[4\]\[6\] _05940_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07150_ _01695_ rvsingle.dp.rf.rf\[6\]\[18\] VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07081_ _01648_ _01998_ _01999_ _01600_ _02001_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_42_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07983_ rvsingle.dp.rf.rf\[23\]\[0\] _01646_ _02903_ VGND VGND VPWR VPWR _02904_
+ sky130_fd_sc_hd__o21ai_1
X_09722_ PC[17] _04554_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__nand2_1
X_06934_ rvsingle.dp.rf.rf\[0\]\[22\] rvsingle.dp.rf.rf\[1\]\[22\] _01562_ VGND VGND
+ VPWR VPWR _01855_ sky130_fd_sc_hd__mux2_1
X_09653_ PC[10] _04475_ PC[11] VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__a21oi_1
X_06865_ _01646_ rvsingle.dp.rf.rf\[31\]\[23\] _01648_ _01785_ VGND VGND VPWR VPWR
+ _01786_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_97_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08604_ rvsingle.dp.rf.rf\[5\]\[12\] VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09584_ _04367_ _04432_ _04437_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[5\] sky130_fd_sc_hd__o21ai_1
X_06796_ _01716_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__buf_4
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08535_ rvsingle.dp.rf.rf\[16\]\[13\] rvsingle.dp.rf.rf\[17\]\[13\] rvsingle.dp.rf.rf\[18\]\[13\]
+ rvsingle.dp.rf.rf\[19\]\[13\] _01416_ _01696_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08466_ rvsingle.dp.rf.rf\[25\]\[9\] _02288_ _01436_ _03386_ VGND VGND VPWR VPWR
+ _03387_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07417_ rvsingle.dp.rf.rf\[3\]\[7\] _01498_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__or2b_1
XFILLER_0_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08397_ _01178_ Instr[29] VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07348_ rvsingle.dp.rf.rf\[13\]\[7\] _01687_ _02268_ VGND VGND VPWR VPWR _02269_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07279_ _01469_ rvsingle.dp.rf.rf\[0\]\[16\] VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09018_ _03930_ _01223_ _01189_ _03937_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10290_ _04719_ _05019_ _05020_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold160 rvsingle.dp.rf.rf\[11\]\[11\] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 rvsingle.dp.rf.rf\[5\]\[21\] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 rvsingle.dp.rf.rf\[4\]\[20\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 rvsingle.dp.rf.rf\[1\]\[4\] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
X_12931_ clknet_leaf_116_clk _00389_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ clknet_leaf_2_clk _00320_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _05867_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__clkbuf_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ clknet_leaf_16_clk _00251_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _04722_ _04723_ _04724_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__or3b_1
XFILLER_0_139_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11675_ _05796_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13414_ clknet_leaf_113_clk _00842_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10626_ _05213_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13345_ clknet_leaf_79_clk rvsingle.dp.PCNext\[22\] _00022_ VGND VGND VPWR VPWR PC[22]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10557_ _05113_ _05114_ _05115_ _05061_ _05173_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__o311a_1
XFILLER_0_51_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13276_ clknet_leaf_129_clk _00734_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10488_ _05131_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__clkbuf_1
X_12227_ _06069_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12158_ _06049_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11109_ _05099_ _05457_ net110 VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__a21oi_1
X_12089_ _04759_ net629 _06010_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__mux2_1
X_06650_ _01559_ rvsingle.dp.rf.rf\[6\]\[21\] VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06581_ _01110_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08320_ rvsingle.dp.rf.rf\[11\]\[8\] _01508_ _02059_ VGND VGND VPWR VPWR _03241_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08251_ _01619_ rvsingle.dp.rf.rf\[10\]\[10\] VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07202_ rvsingle.dp.rf.rf\[23\]\[17\] _01861_ _02122_ VGND VGND VPWR VPWR _02123_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08182_ _03099_ _03100_ _02410_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_132_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07133_ _01493_ rvsingle.dp.rf.rf\[14\]\[18\] _01523_ VGND VGND VPWR VPWR _02054_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07064_ _01973_ _01682_ _01984_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__nand3_4
XFILLER_0_140_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07966_ rvsingle.dp.rf.rf\[29\]\[0\] _01796_ _02485_ VGND VGND VPWR VPWR _02887_
+ sky130_fd_sc_hd__o21ai_1
X_09705_ _04538_ PC[14] _04529_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06917_ _01581_ _01803_ _01837_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__a21oi_2
X_07897_ _02275_ rvsingle.dp.rf.rf\[1\]\[2\] _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_94_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09636_ _04470_ _04471_ _04466_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__or3_1
XFILLER_0_168_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06848_ _01135_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__buf_6
XFILLER_0_168_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09567_ _04139_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__clkbuf_4
X_06779_ _01693_ _01694_ _01698_ _01699_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__a31oi_1
X_08518_ _02395_ _03435_ _03436_ _01502_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_93_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09498_ _04386_ VGND VGND VPWR VPWR WriteData[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08449_ rvsingle.dp.rf.rf\[13\]\[9\] _02288_ _01436_ _03369_ VGND VGND VPWR VPWR
+ _03370_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_93_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11460_ _05364_ _05365_ _05643_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10411_ _04859_ net245 _05082_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__mux2_1
X_11391_ _05641_ _05604_ _05642_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13130_ clknet_leaf_93_clk _00588_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10342_ _05048_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13061_ clknet_leaf_114_clk _00519_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10273_ _04870_ net580 _05001_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__mux2_1
X_12012_ _04721_ _04920_ _05142_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap6 _02260_ VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__buf_1
X_12914_ clknet_leaf_40_clk _00372_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12845_ clknet_leaf_46_clk _00303_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12776_ clknet_leaf_106_clk _00234_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11727_ _05823_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__clkbuf_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11658_ _05713_ net441 _05775_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10609_ _04782_ net479 _05194_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11589_ _05400_ rvsingle.dp.rf.rf\[11\]\[21\] _05729_ VGND VGND VPWR VPWR _05755_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13328_ clknet_leaf_73_clk rvsingle.dp.PCNext\[5\] _00005_ VGND VGND VPWR VPWR PC[5]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13259_ clknet_leaf_100_clk _00717_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07820_ rvsingle.dp.rf.rf\[19\]\[3\] _01124_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__or2b_1
X_07751_ _02669_ _01437_ _01229_ _02671_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_56_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
X_06702_ _01612_ _01615_ _01616_ _01617_ _01622_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__o311ai_2
X_07682_ _01690_ rvsingle.dp.rf.rf\[18\]\[5\] VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09421_ _03311_ _03316_ _04142_ _03312_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__o211a_1
X_06633_ rvsingle.dp.rf.rf\[11\]\[21\] _01509_ _01553_ VGND VGND VPWR VPWR _01554_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09352_ _04262_ _04264_ _04136_ _04267_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__a31oi_4
X_06564_ _01484_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08303_ _01592_ _03194_ _03217_ _01178_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09283_ _04196_ _04198_ _04137_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__nand3_4
X_06495_ _01327_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__buf_6
XFILLER_0_129_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08234_ rvsingle.dp.rf.rf\[8\]\[10\] rvsingle.dp.rf.rf\[9\]\[10\] rvsingle.dp.rf.rf\[10\]\[10\]
+ rvsingle.dp.rf.rf\[11\]\[10\] _02450_ _01708_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08165_ _03078_ _03080_ _03085_ _02491_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_160_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07116_ _01558_ rvsingle.dp.rf.rf\[22\]\[18\] _01880_ VGND VGND VPWR VPWR _02037_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08096_ _03014_ _01502_ _03016_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__nand3_1
XFILLER_0_113_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07047_ _01658_ rvsingle.dp.rf.rf\[20\]\[19\] _01647_ VGND VGND VPWR VPWR _01968_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_100_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08998_ rvsingle.dp.rf.rf\[20\]\[27\] rvsingle.dp.rf.rf\[21\]\[27\] rvsingle.dp.rf.rf\[22\]\[27\]
+ rvsingle.dp.rf.rf\[23\]\[27\] _01337_ _01201_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__mux4_1
X_07949_ rvsingle.dp.rf.rf\[6\]\[0\] _01675_ _01596_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_67_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_16
X_10960_ _05408_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09619_ _04467_ _04453_ _04469_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[8\] sky130_fd_sc_hd__o21ai_1
X_10891_ _05363_ _05315_ _05366_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12630_ clknet_leaf_33_clk _00088_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12561_ clknet_leaf_48_clk _01045_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11512_ _05708_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12492_ clknet_leaf_50_clk _00976_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11443_ _05352_ rvsingle.dp.rf.rf\[13\]\[23\] _05668_ VGND VGND VPWR VPWR _05671_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11374_ _05354_ rvsingle.dp.rf.rf\[14\]\[24\] _05629_ VGND VGND VPWR VPWR _05633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13113_ clknet_leaf_18_clk _00571_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10325_ _05039_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ clknet_leaf_61_clk _00502_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10256_ _04977_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__buf_8
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10187_ _04870_ net748 _04952_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_58_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12828_ clknet_leaf_147_clk _00286_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ clknet_leaf_7_clk _00217_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06280_ _01202_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold704 rvsingle.dp.rf.rf\[1\]\[8\] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 rvsingle.dp.rf.rf\[11\]\[1\] VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold726 rvsingle.dp.rf.rf\[13\]\[8\] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 rvsingle.dp.rf.rf\[31\]\[8\] VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold748 rvsingle.dp.rf.rf\[28\]\[25\] VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ _04786_ net570 _04741_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__mux2_1
Xhold759 rvsingle.dp.rf.rf\[2\]\[25\] VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08921_ _03836_ _03837_ _03838_ _03841_ _03782_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08852_ _01927_ _03772_ _01836_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__o21a_1
X_07803_ rvsingle.dp.rf.rf\[31\]\[3\] _01752_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__or2b_1
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08783_ _01471_ _03701_ _02543_ _03703_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07734_ _01777_ _02651_ _02652_ _01599_ _02654_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__o311ai_2
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07665_ _02583_ _01689_ _01702_ _02585_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09404_ DataAdr[7] DataAdr[10] VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__nor2_1
X_06616_ _01083_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__buf_6
X_07596_ _01614_ rvsingle.dp.rf.rf\[30\]\[4\] VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09335_ _04165_ _02265_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__nand2_2
XFILLER_0_137_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06547_ _01190_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__buf_6
XFILLER_0_118_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09266_ _04179_ _04181_ _04137_ _04183_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_75_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06478_ _01089_ rvsingle.dp.rf.rf\[11\]\[28\] _01261_ _01399_ VGND VGND VPWR VPWR
+ _01400_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08217_ _02093_ _03132_ _03137_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_132_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09197_ _04114_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__nor2_2
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08148_ _03065_ _03066_ _03068_ _01131_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_120_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08079_ rvsingle.dp.rf.rf\[1\]\[1\] _01124_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__or2b_1
X_10110_ net99 VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__inv_2
X_11090_ _05460_ net162 _05178_ _05464_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10041_ _04740_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__buf_6
Xhold20 rvsingle.dp.rf.rf\[3\]\[18\] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 rvsingle.dp.rf.rf\[11\]\[20\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 rvsingle.dp.rf.rf\[27\]\[3\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 rvsingle.dp.rf.rf\[30\]\[0\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 rvsingle.dp.rf.rf\[9\]\[31\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 rvsingle.dp.rf.rf\[25\]\[6\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 rvsingle.dp.rf.rf\[11\]\[3\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 rvsingle.dp.rf.rf\[3\]\[14\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _04852_ net354 _05960_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10943_ _04839_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10874_ _05337_ _05338_ _05339_ _05084_ net319 VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__o41a_1
XFILLER_0_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12613_ clknet_leaf_115_clk _00071_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12544_ clknet_leaf_117_clk _01028_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12475_ clknet_leaf_136_clk _00959_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11426_ _05212_ net720 _05657_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_6 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11357_ _05291_ rvsingle.dp.rf.rf\[14\]\[16\] _05618_ VGND VGND VPWR VPWR _05624_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10308_ _05030_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11288_ _05586_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__clkbuf_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ clknet_leaf_125_clk _00485_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10239_ _04992_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07450_ _02358_ _02370_ _01146_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__nand3_4
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06401_ _01232_ _01318_ _01320_ _01322_ _01224_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07381_ _01444_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__buf_6
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09120_ rvsingle.dp.rf.rf\[19\]\[26\] _03778_ _04039_ VGND VGND VPWR VPWR _04040_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06332_ _01095_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__buf_8
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09051_ _01603_ rvsingle.dp.rf.rf\[12\]\[27\] VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06263_ _01085_ WriteData[30] _01180_ _01185_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__a211o_1
XFILLER_0_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08002_ _01327_ rvsingle.dp.rf.rf\[28\]\[0\] VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06194_ _01117_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold501 rvsingle.dp.rf.rf\[15\]\[9\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold512 rvsingle.dp.rf.rf\[14\]\[26\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 rvsingle.dp.rf.rf\[25\]\[14\] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold534 rvsingle.dp.rf.rf\[29\]\[12\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 rvsingle.dp.rf.rf\[26\]\[5\] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold556 rvsingle.dp.rf.rf\[12\]\[26\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold567 rvsingle.dp.rf.rf\[22\]\[23\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 rvsingle.dp.rf.rf\[8\]\[1\] VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 rvsingle.dp.rf.rf\[20\]\[25\] VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _04772_ _04458_ _04743_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__mux2_8
XFILLER_0_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08904_ _01248_ _03814_ _03824_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__and3_2
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _04422_ _04423_ _04710_ _04711_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _03650_ _03743_ _03729_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__o21ai_1
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _01498_ rvsingle.dp.rf.rf\[2\]\[15\] VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__or2_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ _02634_ _02635_ _02637_ _02323_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__o211ai_1
X_08697_ _02485_ _03614_ _03615_ _02410_ _03617_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__o311ai_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07648_ _02561_ _02568_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__nand2_4
XFILLER_0_95_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07579_ _01878_ rvsingle.dp.rf.rf\[12\]\[4\] VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09318_ _04051_ _04231_ _04232_ _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__o22a_2
XFILLER_0_8_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10590_ _04719_ _05191_ _05192_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09249_ _03770_ _04145_ _04147_ _04167_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_91_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12260_ _05168_ _05847_ _06077_ net128 VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11211_ _05544_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__clkbuf_1
X_12191_ net141 _06049_ _06038_ _05766_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11142_ _05506_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11073_ _04796_ _05145_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__nand2_1
X_10024_ _04425_ _04583_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11975_ _05954_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10926_ _05207_ rvsingle.dp.rf.rf\[18\]\[12\] _05387_ VGND VGND VPWR VPWR _05389_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10857_ _05346_ _05069_ _05068_ _05320_ net39 VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ _04863_ net413 _05298_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__mux2_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12527_ clknet_leaf_39_clk _01011_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12458_ clknet_leaf_82_clk _00942_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11409_ _05381_ net753 _05646_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__mux2_1
X_12389_ clknet_leaf_111_clk _00873_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06950_ _01559_ rvsingle.dp.rf.rf\[30\]\[22\] VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__nor2_1
X_06881_ _01788_ _01801_ _01682_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08620_ rvsingle.dp.rf.rf\[23\]\[12\] _02005_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__and2b_1
X_08551_ _03469_ _01716_ _01460_ _03471_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__a211o_1
X_07502_ _01658_ rvsingle.dp.rf.rf\[6\]\[6\] _01654_ _02422_ VGND VGND VPWR VPWR _02423_
+ sky130_fd_sc_hd__o211ai_1
X_08482_ _01247_ _03397_ _03382_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07433_ rvsingle.dp.rf.rf\[29\]\[7\] _01618_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07364_ _01307_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09103_ _02236_ _04020_ _04022_ _01157_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_72_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06315_ _01232_ _01235_ _01237_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07295_ rvsingle.dp.rf.rf\[17\]\[16\] _01488_ _01497_ _02215_ VGND VGND VPWR VPWR
+ _02216_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_143_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09034_ _01106_ _03951_ _03953_ _02236_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__o211ai_2
X_06246_ Instr[5] VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold320 rvsingle.dp.rf.rf\[26\]\[23\] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold331 rvsingle.dp.rf.rf\[0\]\[28\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ _01100_ rvsingle.dp.rf.rf\[4\]\[30\] VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__or2_1
Xhold342 rvsingle.dp.rf.rf\[1\]\[11\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 rvsingle.dp.rf.rf\[26\]\[11\] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 rvsingle.dp.rf.rf\[18\]\[29\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 rvsingle.dp.rf.rf\[4\]\[24\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold386 rvsingle.dp.rf.rf\[4\]\[16\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 rvsingle.dp.rf.rf\[10\]\[9\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
X_09936_ _04426_ _04757_ _04758_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__a21o_4
XFILLER_0_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _04674_ _04676_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__o21bai_2
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _03647_ _03649_ _03645_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__and3_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _04590_ PC[24] VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__or2_1
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _04833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08749_ rvsingle.dp.rf.rf\[27\]\[15\] _01508_ _03669_ VGND VGND VPWR VPWR _03670_
+ sky130_fd_sc_hd__o21ai_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _05983_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 ReadData[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11760_ _05740_ net649 _05837_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__mux2_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_259 _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10711_ _05259_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _05804_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10642_ _04859_ net567 _05219_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13361_ clknet_leaf_56_clk _00789_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10573_ _04879_ _04881_ _04880_ _05058_ _04876_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__o311a_2
XFILLER_0_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12312_ _04777_ rvsingle.dp.rf.rf\[30\]\[8\] _06099_ VGND VGND VPWR VPWR _06107_
+ sky130_fd_sc_hd__mux2_1
X_13292_ clknet_leaf_93_clk _00750_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12243_ _04746_ net636 _06074_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12174_ _05004_ _05342_ _06052_ net97 VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11125_ _05497_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__clkbuf_1
X_11056_ _05457_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__clkbuf_8
X_10007_ _04817_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__buf_2
XFILLER_0_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11958_ _05945_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10909_ _04765_ rvsingle.dp.rf.rf\[18\]\[5\] _05373_ VGND VGND VPWR VPWR _05379_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11889_ _05496_ rvsingle.dp.rf.rf\[6\]\[6\] _05902_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07080_ _01619_ rvsingle.dp.rf.rf\[2\]\[19\] _01620_ _02000_ VGND VGND VPWR VPWR
+ _02001_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_80_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07982_ rvsingle.dp.rf.rf\[22\]\[0\] _01797_ _01104_ VGND VGND VPWR VPWR _02903_
+ sky130_fd_sc_hd__o21a_1
X_06933_ _01565_ _01850_ _01852_ _01853_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__a31o_1
X_09721_ _04560_ _04562_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06864_ _01125_ rvsingle.dp.rf.rf\[30\]\[23\] VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__or2_1
X_09652_ PC[10] PC[11] _04475_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__and3_1
X_08603_ _03516_ _03518_ _01505_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09583_ _04366_ _04435_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__nand3_1
X_06795_ _01307_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08534_ _03453_ _01084_ _03142_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08465_ _01349_ rvsingle.dp.rf.rf\[24\]\[9\] VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07416_ _01519_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08396_ _03314_ _03316_ _03311_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__o21bai_2
X_07347_ _01306_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__buf_4
XFILLER_0_116_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07278_ rvsingle.dp.rf.rf\[4\]\[16\] rvsingle.dp.rf.rf\[5\]\[16\] rvsingle.dp.rf.rf\[6\]\[16\]
+ rvsingle.dp.rf.rf\[7\]\[16\] _01242_ _01200_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09017_ _02191_ _03931_ _03936_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_104_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06229_ _01152_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold150 rvsingle.dp.rf.rf\[9\]\[3\] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 rvsingle.dp.rf.rf\[8\]\[20\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 rvsingle.dp.rf.rf\[11\]\[14\] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 rvsingle.dp.rf.rf\[17\]\[15\] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold194 rvsingle.dp.rf.rf\[3\]\[12\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
X_09919_ _04121_ _04713_ ReadData[2] _04364_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__a31o_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ clknet_leaf_141_clk _00388_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ clknet_leaf_143_clk _00319_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _05377_ rvsingle.dp.rf.rf\[23\]\[4\] _05863_ VGND VGND VPWR VPWR _05867_
+ sky130_fd_sc_hd__mux2_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ clknet_leaf_31_clk _00250_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _05721_ _05831_ _05833_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__a21oi_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _05724_ rvsingle.dp.rf.rf\[10\]\[1\] _05795_ VGND VGND VPWR VPWR _05796_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13413_ clknet_leaf_112_clk _00841_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10625_ _05212_ rvsingle.dp.rf.rf\[22\]\[15\] _05205_ VGND VGND VPWR VPWR _05213_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10556_ _04827_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13344_ clknet_leaf_78_clk rvsingle.dp.PCNext\[21\] _00021_ VGND VGND VPWR VPWR PC[21]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10487_ _04859_ net528 _05126_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__mux2_1
X_13275_ clknet_leaf_23_clk _00733_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12226_ _06069_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12157_ _06051_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_1
X_11108_ _04721_ _04924_ _05367_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__and3_2
X_12088_ _06013_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__clkbuf_1
X_11039_ _05452_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06580_ rvsingle.dp.rf.rf\[25\]\[21\] _01493_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__or2b_1
XFILLER_0_115_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08250_ _02375_ Instr[30] VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__nand2_2
XFILLER_0_157_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07201_ _01763_ rvsingle.dp.rf.rf\[22\]\[17\] _01777_ VGND VGND VPWR VPWR _02122_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08181_ rvsingle.dp.rf.rf\[15\]\[11\] _01508_ _03101_ VGND VGND VPWR VPWR _03102_
+ sky130_fd_sc_hd__o21ai_2
X_07132_ rvsingle.dp.rf.rf\[13\]\[18\] _01540_ _01543_ VGND VGND VPWR VPWR _02053_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_171_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07063_ _01978_ _01983_ _01116_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07965_ rvsingle.dp.rf.rf\[28\]\[0\] _01126_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__nor2_1
X_09704_ PC[16] _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__xnor2_1
X_06916_ _01591_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__buf_4
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07896_ _01725_ rvsingle.dp.rf.rf\[0\]\[2\] _01454_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09635_ _04483_ PC[8] Instr[28] _04470_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__a31o_1
X_06847_ _01599_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06778_ _01216_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__buf_8
X_09566_ PC[2] PC[3] PC[4] VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__and3_1
X_08517_ _01087_ rvsingle.dp.rf.rf\[13\]\[13\] _03437_ VGND VGND VPWR VPWR _03438_
+ sky130_fd_sc_hd__o21ai_1
X_09497_ _04377_ _03537_ _03560_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__and3_2
XFILLER_0_92_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08448_ _01349_ rvsingle.dp.rf.rf\[12\]\[9\] VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08379_ rvsingle.dp.rf.rf\[25\]\[8\] _01901_ _02285_ _03299_ VGND VGND VPWR VPWR
+ _03300_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10410_ _05086_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11390_ _05364_ _05365_ _05604_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10341_ _04863_ net229 _05044_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13060_ clknet_leaf_123_clk _00518_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10272_ _05010_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12011_ _05971_ _05937_ _05972_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__o21ai_1
X_12913_ clknet_leaf_42_clk _00371_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xmax_cap7 _01069_ VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__buf_2
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ clknet_leaf_51_clk _00302_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ clknet_leaf_98_clk _00233_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _04876_ net550 _05817_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__mux2_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11657_ _05785_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10608_ _05202_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11588_ net31 _05726_ _05754_ _05737_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13327_ clknet_leaf_76_clk rvsingle.dp.PCNext\[4\] _00004_ VGND VGND VPWR VPWR PC[4]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10539_ _04879_ _04881_ _04880_ _05061_ _04785_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__o311a_1
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13258_ clknet_leaf_102_clk _00716_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12209_ _05898_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__inv_2
X_13189_ clknet_leaf_125_clk _00647_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07750_ _02288_ rvsingle.dp.rf.rf\[3\]\[3\] _01433_ _02670_ VGND VGND VPWR VPWR _02671_
+ sky130_fd_sc_hd__o211a_1
X_06701_ _01619_ rvsingle.dp.rf.rf\[14\]\[20\] _01620_ _01621_ VGND VGND VPWR VPWR
+ _01622_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07681_ rvsingle.dp.rf.rf\[17\]\[5\] _02271_ _02268_ _02601_ VGND VGND VPWR VPWR
+ _02602_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06632_ _01137_ rvsingle.dp.rf.rf\[10\]\[21\] _01552_ VGND VGND VPWR VPWR _01553_
+ sky130_fd_sc_hd__o21a_1
X_09420_ _03313_ _03317_ _04153_ _04156_ _04158_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09351_ _04265_ _03454_ _04142_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__o211a_1
X_06563_ _01064_ _01073_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08302_ _01960_ _02102_ _03171_ _03218_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09282_ _04055_ _04193_ _03984_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_118_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06494_ _01411_ _01412_ _01414_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__a21o_1
X_08233_ _03145_ _03147_ _01187_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08164_ _03082_ _01111_ _03084_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__nand3_1
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07115_ rvsingle.dp.rf.rf\[21\]\[18\] _01878_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__and2b_1
XFILLER_0_160_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08095_ rvsingle.dp.rf.rf\[15\]\[1\] _01087_ _03015_ VGND VGND VPWR VPWR _03016_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07046_ _01655_ _01963_ _01964_ _01768_ _01966_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_30_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08997_ _03916_ _01189_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07948_ rvsingle.dp.rf.rf\[5\]\[0\] _01796_ _01092_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o21ai_1
X_07879_ Instr[3] Instr[2] Instr[9] _02799_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__or4_2
XFILLER_0_98_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09618_ _04454_ _04455_ _04468_ _04459_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_168_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10890_ _05364_ _05365_ _05315_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09549_ _04397_ _04367_ _04405_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[2\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12560_ clknet_leaf_68_clk _01044_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11511_ _05300_ rvsingle.dp.rf.rf\[12\]\[22\] _05706_ VGND VGND VPWR VPWR _05708_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12491_ clknet_leaf_64_clk _00975_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11442_ _05670_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11373_ _05632_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10324_ _04818_ net597 _05033_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__mux2_1
X_13112_ clknet_leaf_18_clk _00570_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ net144 _04978_ _05000_ _04985_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__a22o_1
X_13043_ clknet_leaf_26_clk _00501_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10186_ _04956_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12827_ clknet_leaf_142_clk _00285_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ clknet_leaf_34_clk _00216_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11709_ _05439_ net412 _05806_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12689_ clknet_leaf_67_clk _00147_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold705 rvsingle.dp.rf.rf\[29\]\[20\] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 rvsingle.dp.rf.rf\[30\]\[21\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold727 rvsingle.dp.rf.rf\[8\]\[25\] VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 rvsingle.dp.rf.rf\[24\]\[17\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold749 rvsingle.dp.rf.rf\[30\]\[6\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__dlygate4sd3_1
X_08920_ rvsingle.dp.rf.rf\[31\]\[25\] _03839_ _03840_ VGND VGND VPWR VPWR _03841_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08851_ _01838_ _01804_ _01834_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07802_ rvsingle.dp.rf.rf\[29\]\[3\] _01498_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__and2b_1
X_08782_ rvsingle.dp.rf.rf\[29\]\[15\] _02929_ _01307_ _03702_ VGND VGND VPWR VPWR
+ _03703_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07733_ rvsingle.dp.rf.rf\[19\]\[5\] _01087_ _02653_ VGND VGND VPWR VPWR _02654_
+ sky130_fd_sc_hd__o21ai_1
X_07664_ _01687_ rvsingle.dp.rf.rf\[3\]\[5\] _01455_ _02584_ VGND VGND VPWR VPWR _02585_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09403_ _04315_ _04299_ _04316_ VGND VGND VPWR VPWR DataAdr[10] sky130_fd_sc_hd__a21o_4
X_06615_ _01517_ _01535_ _01147_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__nand3_2
XFILLER_0_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07595_ _01853_ _02510_ _02515_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__nand3_1
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06546_ _01208_ _01457_ _01466_ _01218_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__o211ai_1
X_09334_ _02211_ _02263_ _03763_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06477_ _01127_ rvsingle.dp.rf.rf\[10\]\[28\] VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__or2_1
X_09265_ _04182_ _04122_ _04141_ _01288_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_63_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08216_ _02543_ _03134_ _03136_ _01217_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_106_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09196_ _01185_ _04111_ _04113_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__nor3_2
XFILLER_0_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08147_ _02379_ rvsingle.dp.rf.rf\[17\]\[11\] _03067_ VGND VGND VPWR VPWR _03068_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_161_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08078_ rvsingle.dp.rf.rf\[3\]\[1\] _01645_ _01596_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07029_ rvsingle.dp.rf.rf\[4\]\[19\] rvsingle.dp.rf.rf\[5\]\[19\] rvsingle.dp.rf.rf\[6\]\[19\]
+ rvsingle.dp.rf.rf\[7\]\[19\] _01417_ _01301_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10040_ _04845_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__buf_2
Xhold10 rvsingle.dp.rf.rf\[25\]\[17\] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 rvsingle.dp.rf.rf\[3\]\[9\] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 rvsingle.dp.rf.rf\[7\]\[31\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 rvsingle.dp.rf.rf\[6\]\[31\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 rvsingle.dp.rf.rf\[17\]\[6\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 rvsingle.dp.rf.rf\[19\]\[20\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 rvsingle.dp.rf.rf\[11\]\[22\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 rvsingle.dp.rf.rf\[19\]\[12\] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _05962_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__clkbuf_1
Xhold98 rvsingle.dp.rf.rf\[1\]\[14\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
X_10942_ _05397_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10873_ _05355_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12612_ clknet_leaf_107_clk _00070_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12543_ clknet_leaf_1_clk _01027_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12474_ clknet_leaf_5_clk _00958_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11425_ _05661_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11356_ _05623_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10307_ _04778_ net469 _05022_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11287_ _05291_ net803 _05580_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13026_ clknet_leaf_132_clk _00484_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10238_ _04782_ rvsingle.dp.rf.rf\[27\]\[9\] _04989_ VGND VGND VPWR VPWR _04992_
+ sky130_fd_sc_hd__mux2_1
X_10169_ _04947_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06400_ _01202_ _01321_ _01209_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07380_ _02093_ _02294_ _02300_ _01221_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06331_ _01107_ _01253_ _01113_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09050_ _03924_ _01127_ _01106_ _03969_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06262_ _01184_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08001_ rvsingle.dp.rf.rf\[31\]\[0\] _01423_ _01427_ VGND VGND VPWR VPWR _02922_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06193_ _01116_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold502 rvsingle.dp.rf.rf\[31\]\[26\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 rvsingle.dp.rf.rf\[0\]\[12\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 rvsingle.dp.rf.rf\[2\]\[18\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold535 rvsingle.dp.rf.rf\[9\]\[29\] VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 rvsingle.dp.rf.rf\[22\]\[26\] VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 rvsingle.dp.rf.rf\[18\]\[10\] VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold568 rvsingle.dp.rf.rf\[23\]\[24\] VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold579 rvsingle.dp.rf.rf\[6\]\[26\] VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ DataAdr[7] ReadData[7] _04750_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08903_ _01219_ _03817_ _03823_ _01450_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ PC[29] PC[30] PC[31] _04681_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__nand4_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ net820 _03483_ _03565_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__o21ai_4
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ rvsingle.dp.rf.rf\[1\]\[15\] _02478_ _01647_ VGND VGND VPWR VPWR _03686_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _01675_ rvsingle.dp.rf.rf\[28\]\[5\] _02636_ _01667_ VGND VGND VPWR VPWR
+ _02637_ sky130_fd_sc_hd__o211ai_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08696_ _01539_ rvsingle.dp.rf.rf\[21\]\[14\] _03616_ VGND VGND VPWR VPWR _03617_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07647_ _01711_ _02562_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07578_ rvsingle.dp.rf.rf\[15\]\[4\] _01539_ _01520_ VGND VGND VPWR VPWR _02499_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_165_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09317_ _04055_ _04193_ _04136_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06529_ _01187_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__buf_8
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09248_ _04165_ _02101_ _04166_ _03768_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09179_ _01134_ _04094_ _04096_ _04098_ _01157_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__o221a_1
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11210_ _05209_ rvsingle.dp.rf.rf\[29\]\[13\] _05541_ VGND VGND VPWR VPWR _05544_
+ sky130_fd_sc_hd__mux2_1
X_12190_ _04870_ _05766_ _05316_ _06061_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11141_ _05391_ rvsingle.dp.rf.rf\[16\]\[14\] _05499_ VGND VGND VPWR VPWR _05506_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11072_ _05371_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__buf_4
X_10023_ _04751_ _04284_ _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11974_ _04801_ rvsingle.dp.rf.rf\[4\]\[13\] _05949_ VGND VGND VPWR VPWR _05954_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10925_ _05388_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10856_ _04823_ _04726_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10787_ _05302_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12526_ clknet_leaf_72_clk _01010_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12457_ clknet_leaf_96_clk _00941_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11408_ _05652_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12388_ clknet_leaf_122_clk _00872_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11339_ _05614_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13009_ clknet_leaf_57_clk _00467_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06880_ _01791_ _01793_ _01634_ _01800_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08550_ _02929_ rvsingle.dp.rf.rf\[15\]\[13\] _03470_ VGND VGND VPWR VPWR _03471_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07501_ rvsingle.dp.rf.rf\[7\]\[6\] _01557_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__or2b_1
X_08481_ _03400_ _03401_ _01584_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__nand3_2
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07432_ _01862_ rvsingle.dp.rf.rf\[28\]\[7\] VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07363_ _02281_ _01689_ _01702_ _02283_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_128_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09102_ rvsingle.dp.rf.rf\[5\]\[26\] _03839_ _01856_ _04021_ VGND VGND VPWR VPWR
+ _04022_ sky130_fd_sc_hd__o211a_1
X_06314_ _01210_ _01236_ _01224_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07294_ _01595_ rvsingle.dp.rf.rf\[16\]\[16\] VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09033_ _03839_ rvsingle.dp.rf.rf\[27\]\[27\] _03840_ _03952_ VGND VGND VPWR VPWR
+ _03953_ sky130_fd_sc_hd__o211ai_1
X_06245_ _01144_ _01147_ _01154_ _01168_ VGND VGND VPWR VPWR WriteData[30] sky130_fd_sc_hd__o211a_4
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold310 rvsingle.dp.rf.rf\[7\]\[21\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
X_06176_ _01099_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__clkbuf_8
Xhold321 rvsingle.dp.rf.rf\[4\]\[17\] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold332 rvsingle.dp.rf.rf\[19\]\[8\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 rvsingle.dp.rf.rf\[25\]\[16\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold354 rvsingle.dp.rf.rf\[4\]\[22\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 rvsingle.dp.rf.rf\[21\]\[25\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 rvsingle.dp.rf.rf\[2\]\[29\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 rvsingle.dp.rf.rf\[12\]\[16\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 rvsingle.dp.rf.rf\[0\]\[22\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09935_ _04421_ _04424_ _04505_ _04506_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__and4b_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _04671_ _04672_ _04686_ _04687_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__nand4_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _03645_ _03647_ _03649_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__a21oi_1
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _04617_ PC[24] VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__nand2_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _01594_ rvsingle.dp.rf.rf\[26\]\[15\] _01489_ VGND VGND VPWR VPWR _03669_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _04833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_227 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _05983_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 _01097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _01267_ rvsingle.dp.rf.rf\[28\]\[14\] VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _04853_ net670 _05257_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__mux2_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _05428_ net397 _05795_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10641_ _05221_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13360_ clknet_leaf_67_clk _00788_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10572_ net66 _05152_ _05181_ _05157_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12311_ _06106_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13291_ clknet_leaf_100_clk _00749_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12242_ _06075_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12173_ _04802_ _05766_ _05336_ _06056_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11124_ _05496_ rvsingle.dp.rf.rf\[16\]\[6\] _05490_ VGND VGND VPWR VPWR _05497_
+ sky130_fd_sc_hd__mux2_1
X_11055_ _05460_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__clkbuf_8
X_10006_ _04816_ _04556_ _04743_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__mux2_4
XFILLER_0_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11957_ _05534_ net679 _05940_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10908_ _05378_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11888_ _05907_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10839_ _05334_ net342 _05320_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12509_ clknet_leaf_143_clk _00993_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07981_ rvsingle.dp.rf.rf\[21\]\[0\] _01796_ _02485_ _02901_ VGND VGND VPWR VPWR
+ _02902_ sky130_fd_sc_hd__o211ai_1
X_09720_ PC[16] _04546_ _04561_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__a21oi_1
X_06932_ _01155_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__buf_8
X_09651_ _04497_ _04498_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__or2_1
X_06863_ rvsingle.dp.rf.rf\[29\]\[23\] _01646_ _01520_ VGND VGND VPWR VPWR _01784_
+ sky130_fd_sc_hd__o21bai_1
X_08602_ _01620_ _03519_ _03520_ _02323_ _03522_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__o311ai_4
X_09582_ PC[4] _02532_ _04433_ _04434_ _04419_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__a221o_1
X_06794_ rvsingle.dp.rf.rf\[16\]\[20\] rvsingle.dp.rf.rf\[17\]\[20\] _01417_ VGND
+ VGND VPWR VPWR _01715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08533_ _03453_ _01870_ _01485_ _03142_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08464_ rvsingle.dp.rf.rf\[27\]\[9\] _02303_ _03384_ VGND VGND VPWR VPWR _03385_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07415_ _02334_ _02335_ _02329_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08395_ _03315_ _03281_ _01486_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07346_ _01695_ rvsingle.dp.rf.rf\[12\]\[7\] VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07277_ _01222_ _02190_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_61_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09016_ _01461_ _03933_ _03935_ _01447_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06228_ _01151_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06159_ _01082_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__clkbuf_8
Xhold140 rvsingle.dp.rf.rf\[19\]\[4\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 rvsingle.dp.rf.rf\[3\]\[15\] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 rvsingle.dp.rf.rf\[17\]\[22\] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 rvsingle.dp.rf.rf\[19\]\[24\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 rvsingle.dp.rf.rf\[1\]\[12\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 rvsingle.dp.rf.rf\[1\]\[13\] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _04140_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__clkbuf_8
X_09849_ _04422_ _04423_ _04679_ _04427_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ clknet_leaf_148_clk _00318_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _05866_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__clkbuf_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ clknet_leaf_16_clk _00249_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _04973_ _05832_ net79 VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__a21oi_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__buf_6
XFILLER_0_138_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13412_ clknet_leaf_109_clk _00840_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10624_ _04813_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13343_ clknet_leaf_78_clk rvsingle.dp.PCNext\[20\] _00020_ VGND VGND VPWR VPWR PC[20]
+ sky130_fd_sc_hd__dfrtp_4
X_10555_ _05172_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13274_ clknet_leaf_19_clk _00732_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10486_ _05130_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_1
X_12225_ _06069_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12156_ _05728_ net775 _06049_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11107_ _05485_ _05456_ _05486_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__o21ai_1
X_12087_ _04754_ rvsingle.dp.rf.rf\[0\]\[3\] _06010_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__mux2_1
X_11038_ _05266_ net443 _05443_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12989_ clknet_leaf_142_clk _00447_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07200_ rvsingle.dp.rf.rf\[21\]\[17\] _01842_ _01668_ VGND VGND VPWR VPWR _02121_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08180_ _01594_ rvsingle.dp.rf.rf\[14\]\[11\] _01489_ VGND VGND VPWR VPWR _03101_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07131_ _01383_ rvsingle.dp.rf.rf\[12\]\[18\] VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07062_ _01980_ _01632_ _01982_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__nand3_1
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07964_ _01526_ _02867_ _02872_ _02884_ _01593_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09703_ _01226_ _02912_ _01175_ _01171_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__a31o_1
X_06915_ _01804_ _01834_ _01835_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07895_ rvsingle.dp.rf.rf\[3\]\[2\] _02271_ _01300_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09634_ Instr[29] PC[9] VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__or2_1
X_06846_ rvsingle.dp.rf.rf\[1\]\[23\] _01658_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__and2b_1
X_09565_ _04418_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__nor2_1
X_06777_ rvsingle.dp.rf.rf\[15\]\[20\] _01688_ _01697_ VGND VGND VPWR VPWR _01698_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08516_ _01557_ rvsingle.dp.rf.rf\[12\]\[13\] _01103_ VGND VGND VPWR VPWR _03437_
+ sky130_fd_sc_hd__o21ba_1
X_09496_ _03453_ VGND VGND VPWR VPWR WriteData[13] sky130_fd_sc_hd__clkinv_4
XFILLER_0_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08447_ rvsingle.dp.rf.rf\[8\]\[9\] rvsingle.dp.rf.rf\[9\]\[9\] rvsingle.dp.rf.rf\[10\]\[9\]
+ rvsingle.dp.rf.rf\[11\]\[9\] _02176_ _01696_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08378_ _02440_ rvsingle.dp.rf.rf\[24\]\[8\] VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07329_ _01269_ rvsingle.dp.rf.rf\[8\]\[16\] VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10340_ _05047_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10271_ _04863_ net274 _05001_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__mux2_1
X_12010_ _05769_ _05770_ _05937_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12912_ clknet_leaf_52_clk _00370_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12843_ clknet_leaf_88_clk _00301_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ clknet_leaf_113_clk _00232_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _05822_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__clkbuf_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11656_ _05407_ rvsingle.dp.rf.rf\[19\]\[26\] _05775_ VGND VGND VPWR VPWR _05785_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10607_ _04778_ rvsingle.dp.rf.rf\[22\]\[8\] _05194_ VGND VGND VPWR VPWR _05202_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11587_ _04839_ _05732_ _05733_ _05060_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13326_ clknet_leaf_76_clk rvsingle.dp.PCNext\[3\] _00003_ VGND VGND VPWR VPWR PC[3]
+ sky130_fd_sc_hd__dfrtp_4
X_10538_ _05163_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13257_ clknet_leaf_127_clk _00715_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10469_ _05121_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12208_ _05898_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__inv_2
X_13188_ clknet_leaf_137_clk _00646_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_12139_ _05763_ net331 _06031_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__mux2_1
X_06700_ rvsingle.dp.rf.rf\[15\]\[20\] _01255_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__or2b_1
X_07680_ _01690_ rvsingle.dp.rf.rf\[16\]\[5\] VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06631_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__buf_8
X_09350_ _01066_ _01075_ _02261_ _03570_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__a2bb2o_1
X_06562_ Instr[31] VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_48_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08301_ _01246_ _03154_ _03169_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__and3_1
XFILLER_0_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09281_ _04053_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__inv_2
X_06493_ _01348_ _01413_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08232_ _01422_ _03148_ _02438_ _03152_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08163_ rvsingle.dp.rf.rf\[31\]\[11\] _01860_ _03083_ VGND VGND VPWR VPWR _03084_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07114_ _01744_ rvsingle.dp.rf.rf\[20\]\[18\] VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nor2_1
X_08094_ _01096_ rvsingle.dp.rf.rf\[14\]\[1\] _01610_ VGND VGND VPWR VPWR _03015_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07045_ _01256_ rvsingle.dp.rf.rf\[18\]\[19\] _01660_ _01965_ VGND VGND VPWR VPWR
+ _01966_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08996_ _01231_ _03911_ _03915_ _01223_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__o211ai_1
X_07947_ rvsingle.dp.rf.rf\[4\]\[0\] _01643_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07878_ _01068_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09617_ PC[8] _04456_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__xor2_2
X_06829_ rvsingle.dp.rf.rf\[11\]\[23\] _01125_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__or2b_1
XFILLER_0_168_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09548_ _04398_ _04404_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09479_ _04380_ VGND VGND VPWR VPWR WriteData[26] sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_144_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_144_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11510_ _05707_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12490_ clknet_leaf_82_clk _00974_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11441_ _05300_ rvsingle.dp.rf.rf\[13\]\[22\] _05668_ VGND VGND VPWR VPWR _05670_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11372_ _05352_ rvsingle.dp.rf.rf\[14\]\[23\] _05629_ VGND VGND VPWR VPWR _05632_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13111_ clknet_leaf_15_clk _00569_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10323_ _05038_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13042_ clknet_leaf_57_clk _00500_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10254_ _04981_ _04823_ _04982_ _04983_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__and4b_2
X_10185_ _04863_ net742 _04952_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12826_ clknet_leaf_4_clk _00284_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12757_ clknet_leaf_37_clk _00215_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_135_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_135_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _05813_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12688_ clknet_leaf_67_clk _00146_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11639_ _05471_ _05747_ _05779_ net131 VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_4_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold706 rvsingle.dp.rf.rf\[30\]\[4\] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 rvsingle.dp.rf.rf\[15\]\[11\] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold728 rvsingle.dp.rf.rf\[14\]\[27\] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_137_clk _00767_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold739 rvsingle.dp.rf.rf\[20\]\[16\] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08850_ _01589_ _01739_ _03770_ _01840_ _01930_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__a2111o_1
X_07801_ _01642_ rvsingle.dp.rf.rf\[28\]\[3\] VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__nor2_1
X_08781_ _01240_ rvsingle.dp.rf.rf\[28\]\[15\] VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07732_ _01752_ rvsingle.dp.rf.rf\[18\]\[5\] _01610_ VGND VGND VPWR VPWR _02653_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07663_ _01419_ rvsingle.dp.rf.rf\[2\]\[5\] VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__or2_1
X_09402_ _03222_ _03220_ _04142_ _03223_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__o211a_1
X_06614_ _01527_ _01534_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__nand2_1
X_07594_ _02511_ _02512_ _02514_ _01617_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__o211ai_1
X_09333_ _04242_ _04136_ _04243_ _04248_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_165_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06545_ _01458_ _01459_ _01461_ _01465_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_126_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_126_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09264_ _01185_ _01289_ _01347_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06476_ rvsingle.dp.rf.rf\[12\]\[28\] rvsingle.dp.rf.rf\[13\]\[28\] rvsingle.dp.rf.rf\[14\]\[28\]
+ rvsingle.dp.rf.rf\[15\]\[28\] _01099_ _01261_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08215_ _02275_ rvsingle.dp.rf.rf\[27\]\[11\] _01433_ _03135_ VGND VGND VPWR VPWR
+ _03136_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_44_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09195_ _04111_ _04113_ _01185_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08146_ _01779_ rvsingle.dp.rf.rf\[16\]\[11\] _01610_ VGND VGND VPWR VPWR _03067_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08077_ _01847_ rvsingle.dp.rf.rf\[2\]\[1\] VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07028_ _01945_ _01947_ _01208_ _01948_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 rvsingle.dp.rf.rf\[11\]\[7\] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 rvsingle.dp.rf.rf\[1\]\[16\] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 rvsingle.dp.rf.rf\[0\]\[7\] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _01915_ _03893_ _03898_ _01222_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__o211a_1
Xhold44 rvsingle.dp.rf.rf\[23\]\[31\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 rvsingle.dp.rf.rf\[11\]\[31\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 rvsingle.dp.rf.rf\[9\]\[25\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 rvsingle.dp.rf.rf\[24\]\[31\] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _04845_ net278 _05960_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__mux2_1
Xhold88 rvsingle.dp.rf.rf\[9\]\[5\] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 rvsingle.dp.rf.rf\[2\]\[31\] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10941_ _05295_ rvsingle.dp.rf.rf\[18\]\[19\] _05387_ VGND VGND VPWR VPWR _05397_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10872_ _05354_ net244 _05319_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12611_ clknet_leaf_115_clk _00069_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_117_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_117_clk sky130_fd_sc_hd__clkbuf_16
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12542_ clknet_leaf_0_clk _01026_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12473_ clknet_leaf_8_clk _00957_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11424_ _05391_ net697 _05657_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11355_ _05212_ net761 _05618_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10306_ _05029_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__clkbuf_1
X_11286_ _05585_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__clkbuf_1
X_13025_ clknet_leaf_126_clk _00483_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10237_ _04991_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__clkbuf_1
X_10168_ _04818_ rvsingle.dp.rf.rf\[28\]\[16\] _04941_ VGND VGND VPWR VPWR _04947_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10099_ _04426_ _04683_ _04896_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_117_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12809_ clknet_leaf_96_clk _00267_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_108_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_108_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06330_ rvsingle.dp.rf.rf\[2\]\[29\] rvsingle.dp.rf.rf\[3\]\[29\] _01138_ VGND VGND
+ VPWR VPWR _01253_ sky130_fd_sc_hd__mux2_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06261_ _01183_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__buf_4
XFILLER_0_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08000_ _01416_ rvsingle.dp.rf.rf\[30\]\[0\] VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06192_ _01115_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__buf_8
XFILLER_0_53_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold503 rvsingle.dp.rf.rf\[13\]\[29\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 rvsingle.dp.rf.rf\[22\]\[24\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold525 rvsingle.dp.rf.rf\[30\]\[10\] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 rvsingle.dp.rf.rf\[23\]\[19\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold547 rvsingle.dp.rf.rf\[7\]\[20\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _04771_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__clkbuf_1
Xhold558 rvsingle.dp.rf.rf\[22\]\[18\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 rvsingle.dp.rf.rf\[12\]\[21\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ _01703_ _03818_ _03822_ _01478_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ PC[28] PC[29] PC[30] _04663_ PC[31] VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__a41o_1
XFILLER_0_110_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _03746_ _03749_ _03230_ _03753_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__a31oi_2
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _01595_ rvsingle.dp.rf.rf\[0\]\[15\] VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__nor2_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ rvsingle.dp.rf.rf\[29\]\[5\] _01752_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__or2b_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _01267_ rvsingle.dp.rf.rf\[20\]\[14\] _01258_ VGND VGND VPWR VPWR _03616_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07646_ _02564_ _02566_ _02291_ _01446_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07577_ _01780_ rvsingle.dp.rf.rf\[14\]\[4\] VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__nor2_1
X_09316_ _04053_ _04054_ _04193_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06528_ _01230_ _01435_ _01448_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09247_ _02184_ _02265_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06459_ _01095_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__buf_4
XFILLER_0_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09178_ _04097_ _01094_ _01114_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08129_ _02315_ _02982_ _02996_ _01246_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__o211a_2
X_11140_ _05505_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__clkbuf_1
X_11071_ _05470_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10022_ _04140_ _04141_ _04732_ ReadData[19] VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__or4b_1
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11973_ _05953_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10924_ _05334_ net712 _05387_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10855_ _05345_ _05069_ _05068_ _05325_ net22 VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ _04859_ net424 _05298_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__mux2_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ clknet_leaf_44_clk _01009_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12456_ clknet_leaf_106_clk _00940_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11407_ _05496_ net509 _05646_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12387_ clknet_leaf_125_clk _00871_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11338_ _05381_ rvsingle.dp.rf.rf\[14\]\[7\] _05607_ VGND VGND VPWR VPWR _05614_
+ sky130_fd_sc_hd__mux2_1
X_11269_ _05576_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__clkbuf_1
X_13008_ clknet_leaf_55_clk _00466_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07500_ rvsingle.dp.rf.rf\[5\]\[6\] _01613_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__and2b_1
X_08480_ Instr[29] _01083_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__or2_1
X_07431_ _02349_ _02350_ _02351_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07362_ _01695_ rvsingle.dp.rf.rf\[2\]\[7\] _02162_ _02282_ VGND VGND VPWR VPWR _02283_
+ sky130_fd_sc_hd__o211a_1
X_09101_ _01603_ rvsingle.dp.rf.rf\[4\]\[26\] VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06313_ rvsingle.dp.rf.rf\[28\]\[30\] rvsingle.dp.rf.rf\[29\]\[30\] rvsingle.dp.rf.rf\[30\]\[30\]
+ rvsingle.dp.rf.rf\[31\]\[30\] _01196_ _01203_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07293_ rvsingle.dp.rf.rf\[19\]\[16\] _01509_ _01491_ VGND VGND VPWR VPWR _02214_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09032_ _01256_ rvsingle.dp.rf.rf\[26\]\[27\] VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06244_ _01157_ _01160_ _01167_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold300 rvsingle.dp.rf.rf\[1\]\[30\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ _01098_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__clkbuf_8
Xhold311 rvsingle.dp.rf.rf\[17\]\[30\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold322 rvsingle.dp.rf.rf\[27\]\[23\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 rvsingle.dp.rf.rf\[23\]\[16\] VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold344 rvsingle.dp.rf.rf\[20\]\[28\] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold355 rvsingle.dp.rf.rf\[31\]\[7\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 rvsingle.dp.rf.rf\[26\]\[21\] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 rvsingle.dp.rf.rf\[6\]\[29\] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold388 rvsingle.dp.rf.rf\[3\]\[25\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ DataAdr[4] ReadData[4] _04751_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__mux2_1
Xhold399 rvsingle.dp.rf.rf\[16\]\[7\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
X_09865_ PC[30] _01483_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__or2_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ net820 _03483_ _03565_ _03567_ _03572_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_99_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__inv_2
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08747_ rvsingle.dp.rf.rf\[25\]\[15\] _01255_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__and2b_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _04833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _05298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ rvsingle.dp.rf.rf\[31\]\[14\] _01677_ _02320_ VGND VGND VPWR VPWR _03599_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_239 _05983_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _01315_ _02541_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__nand3_2
XFILLER_0_138_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10640_ _04853_ net754 _05219_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10571_ _05113_ _05114_ _05115_ _05061_ _04869_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__o311a_2
XFILLER_0_91_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12310_ _04773_ net622 _06099_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13290_ clknet_leaf_103_clk _00748_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12241_ _04735_ rvsingle.dp.rf.rf\[5\]\[1\] _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12172_ _05337_ _05338_ _05339_ _05003_ net201 VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__o41a_1
XFILLER_0_102_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11123_ _04769_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__buf_2
XFILLER_0_130_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11054_ _05462_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_1
X_10005_ net819 ReadData[16] _04750_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11956_ _05944_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10907_ _05377_ net529 _05373_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__mux2_1
X_11887_ _05534_ net734 _05902_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10838_ _04789_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10769_ _05291_ net739 _05285_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12508_ clknet_leaf_146_clk _00992_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12439_ clknet_leaf_6_clk _00923_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07980_ rvsingle.dp.rf.rf\[20\]\[0\] _01255_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06931_ _01848_ rvsingle.dp.rf.rf\[8\]\[22\] _01851_ _01759_ VGND VGND VPWR VPWR
+ _01852_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09650_ _04481_ _04489_ _04496_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__and3_1
X_06862_ _01643_ rvsingle.dp.rf.rf\[28\]\[23\] VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__nor2_1
X_08601_ _01382_ rvsingle.dp.rf.rf\[14\]\[12\] _01777_ _03521_ VGND VGND VPWR VPWR
+ _03522_ sky130_fd_sc_hd__o211ai_2
X_09581_ _04414_ _04419_ _04433_ _04434_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__o211ai_1
X_06793_ _01701_ _01713_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08532_ _01150_ _01139_ _03429_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_166_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08463_ _02440_ rvsingle.dp.rf.rf\[26\]\[9\] _01243_ VGND VGND VPWR VPWR _03384_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07414_ rvsingle.dp.rf.rf\[1\]\[7\] _01618_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__and2b_1
X_08394_ _01961_ Instr[28] VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07345_ _01931_ _02101_ _02184_ _02265_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__nand4_2
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07276_ _02191_ _02192_ _01222_ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_104_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09015_ _01441_ rvsingle.dp.rf.rf\[3\]\[27\] _01434_ _03934_ VGND VGND VPWR VPWR
+ _03935_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_104_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06227_ _01148_ _01150_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__or2_1
Xhold130 rvsingle.dp.rf.rf\[25\]\[21\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 rvsingle.dp.rf.rf\[3\]\[26\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ Instr[5] _01063_ _01078_ _01067_ _01081_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__o221a_4
Xhold152 rvsingle.dp.rf.rf\[8\]\[9\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 rvsingle.dp.rf.rf\[11\]\[17\] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold174 rvsingle.dp.rf.rf\[3\]\[19\] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 rvsingle.dp.rf.rf\[11\]\[25\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 rvsingle.dp.rf.rf\[19\]\[5\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _04742_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_97_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ PC[28] _04663_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__xor2_1
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _04610_ _04452_ _04615_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[22\] sky130_fd_sc_hd__o21ai_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _05531_ net758 _05863_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__mux2_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ clknet_leaf_31_clk _00248_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11741_ _05830_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__clkbuf_8
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _04738_ _04733_ _05149_ _04739_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__or4b_2
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13411_ clknet_leaf_121_clk _00839_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10623_ _05211_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
X_13342_ clknet_leaf_84_clk rvsingle.dp.PCNext\[19\] _00019_ VGND VGND VPWR VPWR PC[19]
+ sky130_fd_sc_hd__dfrtp_4
X_10554_ _04824_ net478 _05151_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13273_ clknet_leaf_15_clk _00731_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10485_ _04853_ net770 _05126_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__mux2_1
X_12224_ _06069_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__inv_2
X_12155_ _06050_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__clkbuf_1
X_11106_ _05364_ _05365_ _05456_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__o21ai_1
X_12086_ _06012_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_88_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
X_11037_ _05451_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12988_ clknet_leaf_148_clk _00446_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11939_ _05639_ net553 _05924_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_12_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07130_ _01132_ _02048_ _02050_ _01116_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07061_ rvsingle.dp.rf.rf\[31\]\[19\] _01842_ _01981_ VGND VGND VPWR VPWR _01982_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07963_ _01503_ _02875_ _02878_ _01116_ _02883_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__o311ai_4
Xclkbuf_leaf_79_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06914_ _01587_ _01803_ _01066_ _01075_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__a211o_1
X_09702_ _04541_ _04453_ _04545_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[15\] sky130_fd_sc_hd__o21ai_1
X_07894_ _01420_ rvsingle.dp.rf.rf\[2\]\[2\] VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06845_ _01656_ rvsingle.dp.rf.rf\[0\]\[23\] VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09633_ Instr[30] PC[10] VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__or2_1
X_09564_ _04408_ _04417_ _04416_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__a21oi_4
X_06776_ _01695_ rvsingle.dp.rf.rf\[14\]\[20\] _01696_ VGND VGND VPWR VPWR _01697_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08515_ rvsingle.dp.rf.rf\[15\]\[13\] _02627_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__and2b_1
X_09495_ _03644_ VGND VGND VPWR VPWR WriteData[14] sky130_fd_sc_hd__inv_2
XFILLER_0_33_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08446_ _03318_ _03365_ _01486_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08377_ rvsingle.dp.rf.rf\[26\]\[8\] rvsingle.dp.rf.rf\[27\]\[8\] _01707_ VGND VGND
+ VPWR VPWR _03298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07328_ _02245_ _02246_ _02248_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07259_ _02172_ _02174_ _01188_ _02179_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_131_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10270_ _05009_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12911_ clknet_leaf_40_clk _00369_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ clknet_leaf_81_clk _00300_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ clknet_leaf_114_clk _00231_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _05304_ net743 _05817_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__mux2_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11655_ net213 _05778_ _05760_ _05457_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10606_ _05201_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__clkbuf_1
X_11586_ _05167_ _05753_ _05731_ net175 VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10537_ _04782_ net312 _05152_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__mux2_1
X_13325_ clknet_4_12_0_clk rvsingle.dp.PCNext\[2\] _00002_ VGND VGND VPWR VPWR PC[2]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13256_ clknet_leaf_111_clk _00714_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10468_ _04808_ rvsingle.dp.rf.rf\[24\]\[14\] _05110_ VGND VGND VPWR VPWR _05121_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ _05898_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13187_ clknet_leaf_130_clk _00645_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10399_ _05081_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12138_ _06039_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__clkbuf_1
X_12069_ _06002_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_1_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06630_ _01103_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__clkbuf_8
X_06561_ _01481_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08300_ _02469_ _03170_ _03219_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_157_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09280_ _04194_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06492_ _01347_ _01288_ _01290_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08231_ _03149_ _02285_ _01444_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__a211o_1
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08162_ _01544_ rvsingle.dp.rf.rf\[30\]\[11\] _01258_ VGND VGND VPWR VPWR _03083_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07113_ _02028_ _02029_ _01565_ _02033_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_126_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08093_ rvsingle.dp.rf.rf\[13\]\[1\] _01087_ _01667_ _03013_ VGND VGND VPWR VPWR
+ _03014_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_113_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07044_ rvsingle.dp.rf.rf\[19\]\[19\] _01650_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08995_ _03912_ _01310_ _02191_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__a211o_1
X_07946_ _01648_ _02863_ _02864_ _01600_ _02866_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__o311a_1
X_07877_ _01152_ _02774_ _02797_ _01082_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__nand4_4
XFILLER_0_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09616_ _04465_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__xnor2_1
X_06828_ _01745_ _01746_ _01632_ _01748_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06759_ _01092_ _01674_ _01676_ _01679_ _01600_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__o311ai_2
X_09547_ _04400_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09478_ _01962_ _02212_ _04049_ _04031_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_19_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08429_ _01796_ rvsingle.dp.rf.rf\[25\]\[9\] _03349_ VGND VGND VPWR VPWR _03350_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11440_ _05669_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11371_ _05631_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10322_ _04814_ net417 _05033_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__mux2_1
X_13110_ clknet_leaf_25_clk _00568_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13041_ clknet_leaf_57_clk _00499_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10253_ _04999_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__clkbuf_1
X_10184_ _04955_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12825_ clknet_leaf_8_clk _00283_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12756_ clknet_leaf_21_clk _00214_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11707_ _05476_ rvsingle.dp.rf.rf\[10\]\[17\] _05806_ VGND VGND VPWR VPWR _05813_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12687_ clknet_leaf_59_clk _00145_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11638_ _05471_ _05746_ _05779_ net87 VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11569_ _05744_ _05732_ _05733_ _05097_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold707 rvsingle.dp.rf.rf\[28\]\[18\] VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold718 rvsingle.dp.rf.rf\[26\]\[20\] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_14_clk _00766_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold729 rvsingle.dp.rf.rf\[15\]\[19\] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13239_ clknet_leaf_65_clk _00697_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_07800_ _01376_ _02709_ _02720_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__nand3_2
X_08780_ rvsingle.dp.rf.rf\[30\]\[15\] rvsingle.dp.rf.rf\[31\]\[15\] _01903_ VGND
+ VGND VPWR VPWR _03701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07731_ rvsingle.dp.rf.rf\[17\]\[5\] _01566_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07662_ rvsingle.dp.rf.rf\[0\]\[5\] rvsingle.dp.rf.rf\[1\]\[5\] _02176_ VGND VGND
+ VPWR VPWR _02583_ sky130_fd_sc_hd__mux2_1
X_06613_ _01528_ _01529_ _01132_ _01533_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__o211ai_1
X_09401_ _04297_ _04296_ _04135_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07593_ _01513_ rvsingle.dp.rf.rf\[20\]\[4\] _02513_ _02485_ VGND VGND VPWR VPWR
+ _02514_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_75_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06544_ rvsingle.dp.rf.rf\[3\]\[21\] _01296_ _01464_ VGND VGND VPWR VPWR _01465_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09332_ _03907_ _04244_ _03881_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09263_ _04180_ _04059_ _01408_ _01414_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_157_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06475_ _01134_ _01392_ _01394_ _01396_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08214_ _02163_ rvsingle.dp.rf.rf\[26\]\[11\] VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09194_ _04112_ _04110_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08145_ rvsingle.dp.rf.rf\[19\]\[11\] _01860_ _01259_ VGND VGND VPWR VPWR _03066_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08076_ _01188_ _02982_ _02996_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07027_ rvsingle.dp.rf.rf\[12\]\[19\] rvsingle.dp.rf.rf\[13\]\[19\] rvsingle.dp.rf.rf\[14\]\[19\]
+ rvsingle.dp.rf.rf\[15\]\[19\] _01329_ _01456_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__mux4_2
XFILLER_0_113_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold12 rvsingle.dp.rf.rf\[1\]\[18\] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 rvsingle.dp.rf.rf\[24\]\[24\] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _03895_ _01915_ _03897_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__nand3_1
Xhold34 rvsingle.dp.rf.rf\[22\]\[0\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 rvsingle.dp.rf.rf\[5\]\[3\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 rvsingle.dp.rf.rf\[18\]\[31\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 rvsingle.dp.rf.rf\[25\]\[31\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _02849_ _01537_ _01591_ _02798_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__o211ai_4
Xhold78 rvsingle.dp.rf.rf\[9\]\[7\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 rvsingle.dp.rf.rf\[5\]\[7\] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10940_ _05396_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10871_ _04862_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__buf_2
XFILLER_0_168_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12610_ clknet_leaf_128_clk _00068_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12541_ clknet_leaf_143_clk _01025_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12472_ clknet_leaf_34_clk _00956_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11423_ _05660_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11354_ _05622_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__clkbuf_1
X_10305_ _04774_ rvsingle.dp.rf.rf\[26\]\[7\] _05022_ VGND VGND VPWR VPWR _05029_
+ sky130_fd_sc_hd__mux2_1
X_11285_ _05212_ net744 _05580_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__mux2_1
X_13024_ clknet_leaf_118_clk _00482_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10236_ _04778_ net797 _04989_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__mux2_1
X_10167_ _04946_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__clkbuf_1
X_10098_ _04425_ _04895_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12808_ clknet_leaf_123_clk _00266_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12739_ clknet_leaf_116_clk _00197_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06260_ _01064_ _01073_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__nor2_4
XFILLER_0_155_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06191_ Instr[23] VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__buf_12
XFILLER_0_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold504 rvsingle.dp.rf.rf\[28\]\[13\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold515 rvsingle.dp.rf.rf\[28\]\[23\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold526 rvsingle.dp.rf.rf\[6\]\[12\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 rvsingle.dp.rf.rf\[8\]\[16\] VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 rvsingle.dp.rf.rf\[21\]\[20\] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ _04770_ rvsingle.dp.rf.rf\[2\]\[6\] _04741_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__mux2_1
Xhold559 rvsingle.dp.rf.rf\[13\]\[19\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08901_ _03819_ _01437_ _01721_ _03821_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__a211o_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _04704_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ net821 _03141_ _03227_ _03752_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__o22ai_2
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _03675_ _03678_ _02527_ _03683_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07714_ rvsingle.dp.rf.rf\[31\]\[5\] _01860_ _01880_ VGND VGND VPWR VPWR _02635_
+ sky130_fd_sc_hd__o21ai_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ rvsingle.dp.rf.rf\[23\]\[14\] _03258_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__and2b_1
XFILLER_0_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07645_ _01440_ rvsingle.dp.rf.rf\[23\]\[4\] _01696_ _02565_ VGND VGND VPWR VPWR
+ _02566_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07576_ _02493_ _02494_ _02496_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__o21ai_2
X_06527_ _01439_ _01443_ _01445_ _01447_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__a31oi_1
X_09315_ _04230_ _04052_ _04143_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06458_ rvsingle.dp.rf.rf\[28\]\[28\] rvsingle.dp.rf.rf\[29\]\[28\] _01127_ VGND
+ VGND VPWR VPWR _01380_ sky130_fd_sc_hd__mux2_1
X_09246_ _04150_ _04159_ _04164_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09177_ rvsingle.dp.rf.rf\[16\]\[31\] rvsingle.dp.rf.rf\[17\]\[31\] _02212_ VGND
+ VGND VPWR VPWR _04097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06389_ _01310_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__buf_4
XFILLER_0_50_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08128_ _01452_ _02997_ _03047_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08059_ _02976_ _02977_ _02273_ _02979_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__o211ai_1
X_11070_ _05334_ net595 _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__mux2_1
X_10021_ _04829_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__clkbuf_1
X_11972_ _04795_ net680 _05949_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10923_ _05372_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__buf_6
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10854_ _05344_ _04726_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10785_ _05301_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12524_ clknet_leaf_50_clk _01008_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12455_ clknet_leaf_92_clk _00939_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11406_ _05651_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12386_ clknet_leaf_130_clk _00870_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11337_ _05613_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__clkbuf_1
X_11268_ _05381_ net724 _05569_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ clknet_leaf_57_clk _00465_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10219_ _04747_ net639 _04978_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__mux2_1
X_11199_ _05330_ net419 _05528_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07430_ _01599_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__buf_6
XFILLER_0_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07361_ rvsingle.dp.rf.rf\[3\]\[7\] _01828_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09100_ _04018_ _01099_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__a21oi_1
X_06312_ rvsingle.dp.rf.rf\[24\]\[30\] rvsingle.dp.rf.rf\[25\]\[30\] rvsingle.dp.rf.rf\[26\]\[30\]
+ rvsingle.dp.rf.rf\[27\]\[30\] _01225_ _01226_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__mux4_1
X_07292_ _01138_ rvsingle.dp.rf.rf\[18\]\[16\] VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09031_ _03839_ rvsingle.dp.rf.rf\[25\]\[27\] _03950_ VGND VGND VPWR VPWR _03951_
+ sky130_fd_sc_hd__o21ai_1
X_06243_ _01164_ _01166_ _01147_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06174_ _01097_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold301 rvsingle.dp.rf.rf\[28\]\[30\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 rvsingle.dp.rf.rf\[9\]\[9\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold323 rvsingle.dp.rf.rf\[24\]\[30\] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 rvsingle.dp.rf.rf\[9\]\[30\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold345 rvsingle.dp.rf.rf\[21\]\[16\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 rvsingle.dp.rf.rf\[0\]\[8\] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold367 rvsingle.dp.rf.rf\[13\]\[12\] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 rvsingle.dp.rf.rf\[3\]\[24\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _04756_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__clkbuf_1
Xhold389 rvsingle.dp.rf.rf\[25\]\[7\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _01483_ PC[30] VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__nand2_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _03231_ _03406_ _03573_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__nor4_2
XFILLER_0_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _04605_ _04607_ _04619_ _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__or4bb_1
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ _01382_ rvsingle.dp.rf.rf\[24\]\[15\] VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__nor2_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_207 _04884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _05071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _01619_ rvsingle.dp.rf.rf\[30\]\[14\] VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__nor2_1
XANTENNA_229 _05469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _01422_ _02542_ _02548_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07559_ _01619_ rvsingle.dp.rf.rf\[0\]\[4\] VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10570_ _05180_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09229_ _03231_ _03406_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12240_ _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__buf_8
XFILLER_0_161_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12171_ _04796_ _05766_ _05336_ _06055_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11122_ _05495_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__clkbuf_1
X_11053_ _05322_ net654 _05460_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__mux2_1
X_10004_ _04815_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11955_ _04759_ net275 _05940_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10906_ _04759_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__buf_2
XFILLER_0_169_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11886_ _05906_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10837_ _05333_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10768_ _04817_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12507_ clknet_leaf_136_clk _00991_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10699_ _04824_ net630 _05246_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12438_ clknet_leaf_33_clk _00922_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12369_ clknet_leaf_49_clk _00853_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06930_ rvsingle.dp.rf.rf\[9\]\[22\] _01847_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__or2b_1
X_06861_ _01778_ _01781_ _01768_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__o21ai_1
X_08600_ rvsingle.dp.rf.rf\[15\]\[12\] _01566_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__or2b_1
X_06792_ _01703_ _01704_ _01712_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__o21ai_1
X_09580_ Instr[25] _04429_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08531_ _01377_ _03440_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__nand3_4
XFILLER_0_89_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08462_ rvsingle.dp.rf.rf\[28\]\[9\] rvsingle.dp.rf.rf\[29\]\[9\] rvsingle.dp.rf.rf\[30\]\[9\]
+ rvsingle.dp.rf.rf\[31\]\[9\] _01426_ _01433_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07413_ _01753_ rvsingle.dp.rf.rf\[0\]\[7\] _01551_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08393_ _01960_ _02102_ _01084_ _03232_ _03281_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07344_ _02211_ _02264_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__xor2_4
XFILLER_0_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07275_ _01451_ _02193_ _02195_ _01445_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09014_ _01192_ rvsingle.dp.rf.rf\[2\]\[27\] VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06226_ _01149_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold120 rvsingle.dp.rf.rf\[23\]\[0\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlygate4sd3_1
X_06157_ _01080_ _01063_ _01077_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__nand3_2
Xhold131 rvsingle.dp.rf.rf\[19\]\[13\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 rvsingle.dp.rf.rf\[15\]\[0\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 rvsingle.dp.rf.rf\[7\]\[16\] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold164 rvsingle.dp.rf.rf\[5\]\[0\] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 rvsingle.dp.rf.rf\[11\]\[19\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 rvsingle.dp.rf.rf\[9\]\[21\] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 rvsingle.dp.rf.rf\[16\]\[24\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ _04736_ net798 _04741_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _04673_ _04677_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__xnor2_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _04422_ _04423_ _04614_ _04427_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__o211ai_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _03647_ _03649_ _03645_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__nand3_2
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _04720_ _05830_ _04967_ _04968_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__and4_2
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _05721_ _05792_ _05793_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13410_ clknet_leaf_130_clk _00838_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10622_ _04808_ rvsingle.dp.rf.rf\[22\]\[14\] _05205_ VGND VGND VPWR VPWR _05211_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13341_ clknet_leaf_77_clk rvsingle.dp.PCNext\[18\] _00018_ VGND VGND VPWR VPWR PC[18]
+ sky130_fd_sc_hd__dfrtp_4
X_10553_ _05171_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13272_ clknet_leaf_26_clk _00730_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10484_ _05129_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12223_ _06069_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12154_ _05724_ net684 _06049_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11105_ net57 VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__inv_2
X_12085_ _05728_ rvsingle.dp.rf.rf\[0\]\[2\] _06010_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__mux2_1
X_11036_ _05359_ net698 _05443_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12987_ clknet_leaf_141_clk _00445_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11938_ _05933_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__clkbuf_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11869_ _05769_ _05770_ _05860_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07060_ _01642_ rvsingle.dp.rf.rf\[30\]\[19\] _01596_ VGND VGND VPWR VPWR _01981_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07962_ _02879_ _02880_ _02881_ _02882_ _02488_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__o221ai_4
X_09701_ _04454_ _04455_ _04544_ _04459_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__o211ai_1
X_06913_ _01450_ _01820_ _01833_ _01247_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__o211a_2
XFILLER_0_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07893_ _02808_ _02813_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__nand2_4
X_09632_ Instr[30] PC[10] VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__nand2_1
X_06844_ _01762_ _01764_ _01632_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_156_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09563_ _04408_ _04416_ _04417_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__and3_1
X_06775_ _01299_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__buf_6
X_08514_ _01607_ rvsingle.dp.rf.rf\[14\]\[13\] VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09494_ _03697_ VGND VGND VPWR VPWR WriteData[15] sky130_fd_sc_hd__inv_6
XFILLER_0_77_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08445_ _01960_ _02102_ _03318_ _03365_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08376_ _03287_ _03289_ _03296_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07327_ rvsingle.dp.rf.rf\[13\]\[16\] _01488_ _01543_ _02247_ VGND VGND VPWR VPWR
+ _02248_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_73_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07258_ _01230_ _02175_ _02178_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06209_ _01132_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07189_ _01763_ rvsingle.dp.rf.rf\[30\]\[17\] _01777_ VGND VGND VPWR VPWR _02110_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12910_ clknet_leaf_52_clk _00368_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12841_ clknet_leaf_96_clk _00299_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ clknet_leaf_109_clk _00230_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _05821_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__clkbuf_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _05371_ _05759_ _05779_ net173 VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10605_ _04774_ net575 _05194_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__mux2_1
X_11585_ _04834_ _04972_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__nand2_1
X_13324_ clknet_leaf_93_clk _00782_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10536_ _05162_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13255_ clknet_leaf_110_clk _00713_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10467_ _05120_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12206_ _05898_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__inv_2
X_13186_ clknet_leaf_138_clk _00644_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10398_ _04818_ net343 _05071_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12137_ _05713_ net362 _06031_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12068_ _05713_ net814 _05994_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__mux2_1
X_11019_ _05398_ rvsingle.dp.rf.rf\[31\]\[20\] _05431_ VGND VGND VPWR VPWR _05442_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06560_ _01082_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__buf_4
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06491_ _01406_ _01407_ _01375_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08230_ _01294_ rvsingle.dp.rf.rf\[27\]\[10\] _01243_ _03150_ VGND VGND VPWR VPWR
+ _03151_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08161_ _02379_ rvsingle.dp.rf.rf\[29\]\[11\] _03081_ VGND VGND VPWR VPWR _03082_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07112_ rvsingle.dp.rf.rf\[19\]\[18\] _01861_ _02032_ VGND VGND VPWR VPWR _02033_
+ sky130_fd_sc_hd__o21ai_1
X_08092_ _01606_ rvsingle.dp.rf.rf\[12\]\[1\] VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07043_ rvsingle.dp.rf.rf\[17\]\[19\] _01862_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08994_ _01296_ rvsingle.dp.rf.rf\[31\]\[27\] _01200_ _03913_ VGND VGND VPWR VPWR
+ _03914_ sky130_fd_sc_hd__o211a_1
X_07945_ rvsingle.dp.rf.rf\[3\]\[0\] _01842_ _02865_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__o21ai_1
X_07876_ _02785_ _02796_ _01146_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__nand3_4
X_09615_ Instr[28] PC[8] VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__xnor2_1
X_06827_ _01646_ rvsingle.dp.rf.rf\[15\]\[23\] _01105_ _01747_ VGND VGND VPWR VPWR
+ _01748_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_97_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09546_ _04401_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__or2_1
X_06758_ _01677_ rvsingle.dp.rf.rf\[17\]\[20\] _01678_ VGND VGND VPWR VPWR _01679_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09477_ _04379_ VGND VGND VPWR VPWR WriteData[27] sky130_fd_sc_hd__clkbuf_4
X_06689_ Instr[21] VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__buf_4
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08428_ _02005_ rvsingle.dp.rf.rf\[24\]\[9\] _01530_ VGND VGND VPWR VPWR _03349_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08359_ _03261_ _03268_ _01146_ _03279_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_46_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11370_ _05300_ rvsingle.dp.rf.rf\[14\]\[22\] _05629_ VGND VGND VPWR VPWR _05631_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10321_ _05037_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13040_ clknet_leaf_55_clk _00498_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10252_ _04818_ net565 _04989_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__mux2_1
X_10183_ _04859_ net515 _04952_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12824_ clknet_leaf_33_clk _00282_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ clknet_leaf_35_clk _00213_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _05812_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12686_ clknet_leaf_67_clk _00144_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11637_ net189 _05778_ _05745_ _05501_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11568_ _04789_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13307_ clknet_leaf_23_clk _00765_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold708 rvsingle.dp.rf.rf\[14\]\[8\] VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10519_ _04736_ rvsingle.dp.rf.rf\[9\]\[1\] _05152_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__mux2_1
Xhold719 rvsingle.dp.rf.rf\[10\]\[6\] VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11499_ _05701_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13238_ clknet_leaf_62_clk _00696_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13169_ clknet_leaf_58_clk _00627_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07730_ _01650_ rvsingle.dp.rf.rf\[16\]\[5\] VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07661_ _02579_ _01444_ _02581_ _01215_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09400_ _04312_ _04313_ _04314_ _04143_ VGND VGND VPWR VPWR DataAdr[7] sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_133_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06612_ rvsingle.dp.rf.rf\[19\]\[21\] _01488_ _01532_ VGND VGND VPWR VPWR _01533_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07592_ rvsingle.dp.rf.rf\[21\]\[4\] _01267_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09331_ _04246_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__buf_4
X_06543_ _01463_ rvsingle.dp.rf.rf\[2\]\[21\] _01199_ VGND VGND VPWR VPWR _01464_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09262_ _01411_ _01412_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__and2_2
XFILLER_0_7_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06474_ _01395_ _01094_ _01113_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08213_ rvsingle.dp.rf.rf\[25\]\[11\] _01827_ _01308_ _03133_ VGND VGND VPWR VPWR
+ _03134_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_106_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09193_ _01248_ _04076_ _04087_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08144_ _01382_ rvsingle.dp.rf.rf\[18\]\[11\] VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08075_ _02986_ _02988_ _01187_ _02995_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07026_ _01946_ _01717_ _01445_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold13 rvsingle.dp.rf.rf\[1\]\[5\] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ rvsingle.dp.rf.rf\[15\]\[25\] _01297_ _03896_ VGND VGND VPWR VPWR _03897_
+ sky130_fd_sc_hd__o21ai_1
Xhold24 rvsingle.dp.rf.rf\[28\]\[0\] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 rvsingle.dp.rf.rf\[2\]\[0\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 rvsingle.dp.rf.rf\[16\]\[31\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 rvsingle.dp.rf.rf\[17\]\[31\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _01113_ net825 _02800_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__o21ai_2
Xhold68 rvsingle.dp.rf.rf\[27\]\[31\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 rvsingle.dp.rf.rf\[7\]\[0\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _01097_ rvsingle.dp.rf.rf\[24\]\[2\] VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10870_ _05353_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09529_ _04256_ VGND VGND VPWR VPWR DataAdr[17] sky130_fd_sc_hd__clkinv_4
XFILLER_0_94_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12540_ clknet_leaf_151_clk _01024_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12471_ clknet_leaf_6_clk _00955_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11422_ _04801_ net488 _05657_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11353_ _05391_ net604 _05618_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10304_ _05028_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__clkbuf_1
X_11284_ _05584_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13023_ clknet_leaf_13_clk _00481_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10235_ _04990_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__clkbuf_1
X_10166_ _04814_ rvsingle.dp.rf.rf\[28\]\[15\] _04941_ VGND VGND VPWR VPWR _04946_
+ sky130_fd_sc_hd__mux2_1
X_10097_ _04751_ _04184_ _04894_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12807_ clknet_leaf_98_clk _00265_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10999_ _05418_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__buf_6
XFILLER_0_57_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ clknet_leaf_129_clk _00196_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12669_ clknet_leaf_143_clk _00127_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06190_ _01113_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__buf_4
XFILLER_0_114_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold505 rvsingle.dp.rf.rf\[23\]\[20\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold516 rvsingle.dp.rf.rf\[10\]\[10\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 rvsingle.dp.rf.rf\[8\]\[22\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 rvsingle.dp.rf.rf\[2\]\[9\] VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold549 rvsingle.dp.rf.rf\[4\]\[7\] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08900_ _02288_ rvsingle.dp.rf.rf\[15\]\[24\] _01433_ _03820_ VGND VGND VPWR VPWR
+ _03821_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _04701_ _04705_ _04706_ _04707_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__o22ai_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _02469_ _03228_ _03112_ _03751_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__a2bb2oi_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _03679_ _03680_ _01511_ _03682_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__o211ai_2
X_07713_ _01862_ rvsingle.dp.rf.rf\[30\]\[5\] VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08693_ _01763_ rvsingle.dp.rf.rf\[22\]\[14\] VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07644_ _01419_ rvsingle.dp.rf.rf\[22\]\[4\] VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07575_ _02481_ rvsingle.dp.rf.rf\[9\]\[4\] _02495_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09314_ _04002_ _04013_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__nor2_1
X_06526_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09245_ _04161_ _04149_ _04163_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__a21oi_1
X_06457_ rvsingle.dp.rf.rf\[24\]\[28\] rvsingle.dp.rf.rf\[25\]\[28\] rvsingle.dp.rf.rf\[26\]\[28\]
+ rvsingle.dp.rf.rf\[27\]\[28\] _01099_ _01261_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09176_ _01090_ rvsingle.dp.rf.rf\[19\]\[31\] _01120_ _04095_ VGND VGND VPWR VPWR
+ _04096_ sky130_fd_sc_hd__o211a_1
X_06388_ _01309_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08127_ _01065_ _01074_ _03043_ _03046_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08058_ rvsingle.dp.rf.rf\[7\]\[1\] _01295_ _02978_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07009_ _01927_ _01929_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10020_ _04828_ net524 _04791_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11971_ _05952_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__clkbuf_1
X_10922_ _05386_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10853_ _04817_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10784_ _05300_ net463 _05298_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ clknet_leaf_86_clk _01007_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12454_ clknet_leaf_108_clk _00938_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11405_ _05534_ rvsingle.dp.rf.rf\[13\]\[5\] _05646_ VGND VGND VPWR VPWR _05651_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12385_ clknet_leaf_125_clk _00869_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11336_ _05496_ net410 _05607_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__mux2_1
X_11267_ _05575_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13006_ clknet_leaf_55_clk _00464_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10218_ _04979_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11198_ _05537_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__clkbuf_1
X_10149_ _04774_ net809 _04930_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07360_ rvsingle.dp.rf.rf\[0\]\[7\] rvsingle.dp.rf.rf\[1\]\[7\] _01241_ VGND VGND
+ VPWR VPWR _02281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06311_ _01232_ _01233_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07291_ _01128_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__buf_6
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09030_ _01256_ rvsingle.dp.rf.rf\[24\]\[27\] VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06242_ _01114_ _01165_ _01118_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06173_ _01096_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__buf_6
Xhold302 rvsingle.dp.rf.rf\[29\]\[30\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold313 rvsingle.dp.rf.rf\[3\]\[30\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 rvsingle.dp.rf.rf\[3\]\[28\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold335 rvsingle.dp.rf.rf\[16\]\[25\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 rvsingle.dp.rf.rf\[10\]\[16\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 rvsingle.dp.rf.rf\[8\]\[17\] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _04755_ rvsingle.dp.rf.rf\[2\]\[3\] _04741_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__mux2_1
Xhold368 rvsingle.dp.rf.rf\[12\]\[14\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold379 rvsingle.dp.rf.rf\[10\]\[27\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ PC[29] PC[30] _04681_ _04691_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__a31o_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _03648_ _03650_ _03729_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__nand4_2
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _04588_ _04625_ _04609_ _04626_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__or4_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _03662_ _03663_ _03665_ _02488_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _04892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _03588_ _03590_ _02315_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__o211ai_4
XANTENNA_219 _05085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _02543_ _02545_ _02547_ _01446_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__a31oi_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07558_ rvsingle.dp.rf.rf\[3\]\[4\] _02478_ _01523_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06509_ _01421_ _01309_ _01422_ _01429_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07489_ _01110_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__clkbuf_8
X_09228_ _04146_ _01590_ _01739_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__or3b_1
XFILLER_0_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09159_ _04077_ _04078_ _01232_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12170_ _05337_ _05338_ _05339_ _05004_ net194 VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__o41a_1
X_11121_ _04765_ rvsingle.dp.rf.rf\[16\]\[5\] _05490_ VGND VGND VPWR VPWR _05495_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11052_ _05461_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
X_10003_ _04814_ net227 _04791_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11954_ _05943_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10905_ _05376_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11885_ _04759_ net542 _05902_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10836_ _04786_ net489 _05320_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10767_ _05290_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12506_ clknet_leaf_4_clk _00990_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10698_ _05252_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__clkbuf_1
X_12437_ clknet_leaf_36_clk _00921_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12368_ clknet_leaf_72_clk _00852_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11319_ _05364_ _05365_ _05566_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12299_ _06100_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06860_ rvsingle.dp.rf.rf\[25\]\[23\] _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__and2b_1
X_06791_ _01706_ _01710_ _01711_ _01221_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08530_ _01156_ _03445_ _03450_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__nand3_1
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08461_ _01315_ _03374_ _03381_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__nand3_2
XFILLER_0_148_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07412_ _02326_ _02332_ _01505_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__nand3_1
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08392_ _03283_ _03311_ _03312_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__nand3_4
XFILLER_0_147_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07343_ _02258_ _02261_ _02263_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07274_ rvsingle.dp.rf.rf\[25\]\[16\] _01424_ _01716_ _02194_ VGND VGND VPWR VPWR
+ _02195_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09013_ rvsingle.dp.rf.rf\[1\]\[27\] _01441_ _01437_ _03932_ VGND VGND VPWR VPWR
+ _03933_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06225_ _01145_ Instr[21] Instr[22] _01115_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold110 rvsingle.dp.rf.rf\[16\]\[0\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ Instr[1] Instr[0] _01076_ _01079_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__nand4_4
Xhold121 rvsingle.dp.rf.rf\[17\]\[3\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 rvsingle.dp.rf.rf\[1\]\[15\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold143 rvsingle.dp.rf.rf\[11\]\[12\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold154 rvsingle.dp.rf.rf\[27\]\[21\] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 rvsingle.dp.rf.rf\[7\]\[13\] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold176 rvsingle.dp.rf.rf\[3\]\[16\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold187 rvsingle.dp.rf.rf\[10\]\[0\] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 rvsingle.dp.rf.rf\[17\]\[4\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _04740_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__buf_8
XFILLER_0_10_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09846_ _04674_ _04676_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__nor2_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _04612_ _04613_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__nor2_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _01296_ rvsingle.dp.rf.rf\[27\]\[22\] _01434_ _01909_ VGND VGND VPWR VPWR
+ _01910_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _01338_ _01245_ _01201_ _03597_ _03586_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__o311a_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08659_ rvsingle.dp.rf.rf\[0\]\[14\] rvsingle.dp.rf.rf\[1\]\[14\] rvsingle.dp.rf.rf\[2\]\[14\]
+ rvsingle.dp.rf.rf\[3\]\[14\] _01730_ _01433_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__mux4_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11670_ net187 _05792_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10621_ _05210_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13340_ clknet_leaf_77_clk rvsingle.dp.PCNext\[17\] _00017_ VGND VGND VPWR VPWR PC[17]
+ sky130_fd_sc_hd__dfrtp_4
X_10552_ _04818_ net664 _05151_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13271_ clknet_leaf_60_clk _00729_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10483_ _04846_ net436 _05126_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12222_ reset VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12153_ _06048_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__buf_8
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11104_ _05484_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__clkbuf_1
X_12084_ _06011_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__clkbuf_1
X_11035_ _05450_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12986_ clknet_leaf_1_clk _00444_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11937_ _05716_ net377 _05924_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__mux2_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11868_ net44 VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10819_ _05323_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11799_ _05769_ _05770_ _05831_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07961_ rvsingle.dp.rf.rf\[13\]\[0\] _01487_ _01496_ VGND VGND VPWR VPWR _02882_
+ sky130_fd_sc_hd__o21ai_2
X_09700_ _04542_ _04543_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__nor2_1
X_06912_ _01822_ _01824_ _01188_ _01832_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__o211ai_1
X_07892_ _02809_ _02810_ _02543_ _02812_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09631_ _04479_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__inv_2
X_06843_ rvsingle.dp.rf.rf\[5\]\[23\] _01763_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__and2b_1
X_09562_ PC[3] _02748_ _04401_ _04410_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__o22ai_4
X_06774_ _01349_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__buf_8
X_08513_ _03430_ _03431_ _03433_ _01131_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__o211ai_1
X_09493_ _02257_ VGND VGND VPWR VPWR WriteData[16] sky130_fd_sc_hd__inv_4
XFILLER_0_66_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08444_ _03341_ _01481_ _01592_ _03364_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__nand4_2
XFILLER_0_148_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08375_ _02093_ _03290_ _03295_ _01447_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07326_ _01499_ rvsingle.dp.rf.rf\[12\]\[16\] VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07257_ _02093_ _02177_ _01699_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06208_ _01131_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07188_ rvsingle.dp.rf.rf\[29\]\[17\] _01842_ _01668_ VGND VGND VPWR VPWR _02109_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06139_ Instr[1] Instr[0] _01061_ _01062_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__nand4_4
XFILLER_0_112_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09829_ _04422_ _04423_ _04661_ _04427_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__o211ai_1
X_12840_ clknet_leaf_104_clk _00298_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ clknet_leaf_116_clk _00229_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_147_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_147_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _05354_ net259 _05817_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _05784_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _05200_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11584_ _05752_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13323_ clknet_leaf_127_clk _00781_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10535_ _04778_ rvsingle.dp.rf.rf\[9\]\[8\] _05152_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13254_ clknet_leaf_101_clk _00712_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10466_ _04802_ rvsingle.dp.rf.rf\[24\]\[13\] _05110_ VGND VGND VPWR VPWR _05120_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12205_ _05898_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__inv_2
X_13185_ clknet_leaf_133_clk _00643_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10397_ _05080_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__clkbuf_1
X_12136_ _06038_ _05060_ _04924_ _06010_ net180 VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__a32o_1
X_12067_ _06001_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__clkbuf_1
X_11018_ _05441_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_138_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12969_ clknet_leaf_97_clk _00427_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06490_ _01375_ _01406_ _01407_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__nand3_1
XFILLER_0_129_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08160_ _01779_ rvsingle.dp.rf.rf\[28\]\[11\] _01610_ VGND VGND VPWR VPWR _03081_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07111_ _02030_ rvsingle.dp.rf.rf\[18\]\[18\] _02031_ VGND VGND VPWR VPWR _02032_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08091_ _03008_ _03009_ _03010_ _03011_ _01564_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07042_ _01656_ rvsingle.dp.rf.rf\[16\]\[19\] VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08993_ _01432_ rvsingle.dp.rf.rf\[30\]\[27\] VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07944_ rvsingle.dp.rf.rf\[2\]\[0\] _01753_ _01596_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__o21a_1
X_07875_ _01156_ _02790_ _02795_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__nand3_1
X_06826_ _01125_ rvsingle.dp.rf.rf\[14\]\[23\] VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__or2_1
X_09614_ _04462_ _04464_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09545_ _04397_ _02801_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__nor2_1
X_06757_ _01602_ rvsingle.dp.rf.rf\[16\]\[20\] _01551_ VGND VGND VPWR VPWR _01678_
+ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_129_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_129_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09476_ _01154_ _03956_ _03977_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__and3_2
XFILLER_0_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06688_ _01603_ rvsingle.dp.rf.rf\[10\]\[20\] _01605_ _01608_ VGND VGND VPWR VPWR
+ _01609_ sky130_fd_sc_hd__o211a_1
X_08427_ rvsingle.dp.rf.rf\[27\]\[9\] _01796_ _03347_ VGND VGND VPWR VPWR _03348_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08358_ _01853_ _03273_ _03278_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__nand3_1
XFILLER_0_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07309_ _01493_ rvsingle.dp.rf.rf\[30\]\[16\] _01523_ VGND VGND VPWR VPWR _02230_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08289_ _01614_ rvsingle.dp.rf.rf\[26\]\[10\] _02320_ _03209_ VGND VGND VPWR VPWR
+ _03210_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10320_ _04808_ net457 _05033_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10251_ _04998_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_898 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10182_ _04954_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12823_ clknet_leaf_6_clk _00281_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ clknet_leaf_40_clk _00212_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _05344_ net346 _05806_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__mux2_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12685_ clknet_leaf_45_clk _00143_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11636_ net18 _05778_ _05743_ _05501_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11567_ net93 _05726_ _05743_ _05737_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10518_ _05151_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__buf_8
X_13306_ clknet_leaf_19_clk _00764_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold709 rvsingle.dp.rf.rf\[31\]\[6\] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11498_ _05291_ net387 _05695_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13237_ clknet_leaf_10_clk _00695_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10449_ _05109_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13168_ clknet_leaf_71_clk _00626_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12119_ _06029_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__clkbuf_1
X_13099_ clknet_leaf_88_clk _00557_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07660_ rvsingle.dp.rf.rf\[7\]\[5\] _01440_ _02580_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__o21ai_1
X_06611_ _01256_ rvsingle.dp.rf.rf\[18\]\[21\] _01531_ VGND VGND VPWR VPWR _01532_
+ sky130_fd_sc_hd__o21a_1
X_07591_ rvsingle.dp.rf.rf\[23\]\[4\] _02481_ _02320_ VGND VGND VPWR VPWR _02512_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09330_ _04245_ _04122_ _02259_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__or3b_1
X_06542_ _01462_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09261_ _01409_ _04178_ _01414_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__o21bai_2
X_06473_ rvsingle.dp.rf.rf\[0\]\[28\] rvsingle.dp.rf.rf\[1\]\[28\] _01127_ VGND VGND
+ VPWR VPWR _01395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08212_ _02163_ rvsingle.dp.rf.rf\[24\]\[11\] VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09192_ _01248_ _04076_ _04087_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__and4_1
XFILLER_0_117_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08143_ _02668_ _03054_ _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_16_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08074_ _02302_ _02989_ _02994_ _02438_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_114_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07025_ rvsingle.dp.rf.rf\[8\]\[19\] rvsingle.dp.rf.rf\[9\]\[19\] _01469_ VGND VGND
+ VPWR VPWR _01946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold14 rvsingle.dp.rf.rf\[11\]\[9\] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _01193_ rvsingle.dp.rf.rf\[14\]\[25\] _01200_ VGND VGND VPWR VPWR _03896_
+ sky130_fd_sc_hd__o21a_1
Xhold25 rvsingle.dp.rf.rf\[30\]\[31\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 rvsingle.dp.rf.rf\[7\]\[4\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 rvsingle.dp.rf.rf\[20\]\[31\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 rvsingle.dp.rf.rf\[21\]\[31\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _01246_ _02826_ _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__and3_2
Xhold69 rvsingle.dp.rf.rf\[7\]\[15\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
X_07858_ _02775_ _02776_ _02410_ _02778_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__o211ai_1
X_06809_ _01425_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__clkbuf_8
X_07789_ _02005_ rvsingle.dp.rf.rf\[0\]\[3\] VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09528_ _04228_ _04396_ VGND VGND VPWR VPWR DataAdr[15] sky130_fd_sc_hd__nand2_8
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09459_ _04139_ _04363_ _04365_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12470_ clknet_leaf_31_clk _00954_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11421_ _05659_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11352_ _05621_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__clkbuf_1
X_10303_ _04770_ net789 _05022_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11283_ _05391_ rvsingle.dp.rf.rf\[15\]\[14\] _05580_ VGND VGND VPWR VPWR _05584_
+ sky130_fd_sc_hd__mux2_1
X_13022_ clknet_leaf_134_clk _00480_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10234_ _04774_ rvsingle.dp.rf.rf\[27\]\[7\] _04989_ VGND VGND VPWR VPWR _04990_
+ sky130_fd_sc_hd__mux2_1
X_10165_ _04945_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10096_ _04140_ _04141_ _04732_ ReadData[29] VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__or4b_1
XFILLER_0_89_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12806_ clknet_leaf_113_clk _00264_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10998_ _05430_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12737_ clknet_leaf_141_clk _00195_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12668_ clknet_leaf_151_clk _00126_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_955 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11619_ _05721_ _05772_ _05773_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12599_ clknet_leaf_7_clk _00057_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold506 rvsingle.dp.rf.rf\[30\]\[12\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold517 rvsingle.dp.rf.rf\[20\]\[27\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold528 rvsingle.dp.rf.rf\[24\]\[23\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 rvsingle.dp.rf.rf\[24\]\[18\] VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _01482_ _01171_ _01584_ _03750_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ rvsingle.dp.rf.rf\[13\]\[15\] _01487_ _02395_ _03681_ VGND VGND VPWR VPWR
+ _03682_ sky130_fd_sc_hd__o211ai_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _01377_ _02620_ _02632_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__nand3_4
X_08692_ _01531_ _03609_ _03610_ _01131_ _03612_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07643_ rvsingle.dp.rf.rf\[21\]\[4\] _01827_ _01308_ _02563_ VGND VGND VPWR VPWR
+ _02564_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_95_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07574_ _01561_ rvsingle.dp.rf.rf\[8\]\[4\] _01489_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_119_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09313_ _03731_ _04123_ _04211_ _04219_ _04228_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__o311a_1
XFILLER_0_119_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06525_ _01215_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__buf_6
XFILLER_0_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_60_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
X_09244_ _03735_ _04162_ _03756_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06456_ _01377_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__buf_8
XFILLER_0_134_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09175_ _02212_ rvsingle.dp.rf.rf\[18\]\[31\] VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06387_ _01308_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__buf_6
XFILLER_0_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08126_ _03043_ _03046_ _01485_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_32_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08057_ _01468_ rvsingle.dp.rf.rf\[6\]\[1\] _01198_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__o21a_1
X_07008_ _01928_ _01898_ _01925_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08959_ _01085_ WriteData[25] VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__nand2_1
X_11970_ _05744_ net576 _05949_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10921_ _05385_ net557 _05373_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__mux2_1
X_10852_ _05085_ _05343_ _05325_ net132 VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__a2bb2o_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10783_ _04852_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__buf_2
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ clknet_leaf_83_clk _01006_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12453_ clknet_leaf_114_clk _00937_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11404_ _05650_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__clkbuf_1
X_12384_ clknet_leaf_119_clk _00868_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11335_ _05612_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11266_ _05496_ net646 _05569_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__mux2_1
X_10217_ _04736_ net350 _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__mux2_1
X_13005_ clknet_leaf_45_clk _00463_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11197_ _05381_ net444 _05528_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10148_ _04936_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__clkbuf_1
X_10079_ _02909_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_42_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
X_06310_ rvsingle.dp.rf.rf\[16\]\[30\] rvsingle.dp.rf.rf\[17\]\[30\] rvsingle.dp.rf.rf\[18\]\[30\]
+ rvsingle.dp.rf.rf\[19\]\[30\] _01225_ _01226_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07290_ _01317_ _02198_ _02210_ _01248_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06241_ rvsingle.dp.rf.rf\[24\]\[30\] rvsingle.dp.rf.rf\[25\]\[30\] rvsingle.dp.rf.rf\[26\]\[30\]
+ rvsingle.dp.rf.rf\[27\]\[30\] _01128_ _01107_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06172_ _01095_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold303 rvsingle.dp.rf.rf\[5\]\[24\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 rvsingle.dp.rf.rf\[4\]\[8\] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold325 rvsingle.dp.rf.rf\[21\]\[9\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold336 rvsingle.dp.rf.rf\[6\]\[11\] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 rvsingle.dp.rf.rf\[22\]\[21\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold358 rvsingle.dp.rf.rf\[8\]\[28\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__buf_2
Xhold369 rvsingle.dp.rf.rf\[22\]\[17\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ PC[28] PC[29] _04663_ PC[30] VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__a31oi_2
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _03731_ _03732_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__o21ai_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _04549_ _04551_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _01499_ rvsingle.dp.rf.rf\[28\]\[15\] _03664_ _01496_ VGND VGND VPWR VPWR
+ _03665_ sky130_fd_sc_hd__o211ai_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _04978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08675_ _01711_ _03591_ _03595_ _01221_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__o211ai_2
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07626_ rvsingle.dp.rf.rf\[1\]\[4\] _02271_ _02268_ _02546_ VGND VGND VPWR VPWR _02547_
+ sky130_fd_sc_hd__o211ai_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07557_ _01086_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_33_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
X_06508_ _01424_ rvsingle.dp.rf.rf\[31\]\[21\] _01428_ VGND VGND VPWR VPWR _01429_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07488_ rvsingle.dp.rf.rf\[13\]\[6\] _02379_ _01542_ VGND VGND VPWR VPWR _02409_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06439_ _01219_ _01354_ _01360_ _01317_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__a211o_1
X_09227_ _01740_ _01685_ _01737_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_91_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09158_ rvsingle.dp.rf.rf\[20\]\[31\] rvsingle.dp.rf.rf\[21\]\[31\] rvsingle.dp.rf.rf\[22\]\[31\]
+ rvsingle.dp.rf.rf\[23\]\[31\] _01225_ _01226_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08109_ _02364_ _03024_ _03029_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__nand3_1
X_09089_ rvsingle.dp.rf.rf\[16\]\[26\] rvsingle.dp.rf.rf\[17\]\[26\] rvsingle.dp.rf.rf\[18\]\[26\]
+ rvsingle.dp.rf.rf\[19\]\[26\] _01337_ _01302_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__mux4_1
X_11120_ _05494_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__clkbuf_1
X_11051_ _05318_ net471 _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__mux2_1
X_10002_ _04813_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11953_ _05531_ rvsingle.dp.rf.rf\[4\]\[3\] _05940_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10904_ _04755_ rvsingle.dp.rf.rf\[18\]\[3\] _05373_ VGND VGND VPWR VPWR _05376_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11884_ _05905_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10835_ _05332_ _05069_ _05068_ _05325_ net3 VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10766_ _05212_ rvsingle.dp.rf.rf\[20\]\[15\] _05285_ VGND VGND VPWR VPWR _05290_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12505_ clknet_leaf_7_clk _00989_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10697_ _04818_ net345 _05246_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12436_ clknet_leaf_21_clk _00920_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12367_ clknet_leaf_57_clk _00851_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11318_ net70 VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__inv_2
X_12298_ _04735_ rvsingle.dp.rf.rf\[30\]\[1\] _06099_ VGND VGND VPWR VPWR _06100_
+ sky130_fd_sc_hd__mux2_1
X_11249_ _05563_ _05525_ _05564_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06790_ _01444_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__buf_8
X_08460_ _01711_ _03375_ _03380_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07411_ _01523_ _02327_ _02328_ _02329_ _02331_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_147_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08391_ _01960_ _02102_ _01084_ _03232_ _03281_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07342_ _01066_ _01075_ _01587_ _02262_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__o211a_2
XFILLER_0_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07273_ _02176_ rvsingle.dp.rf.rf\[24\]\[16\] VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09012_ _01192_ rvsingle.dp.rf.rf\[0\]\[27\] VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06224_ _01096_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__buf_6
XFILLER_0_170_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold100 rvsingle.dp.rf.rf\[3\]\[5\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06155_ Instr[6] Instr[3] Instr[2] VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__and3_2
XFILLER_0_79_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold111 rvsingle.dp.rf.rf\[6\]\[0\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold122 rvsingle.dp.rf.rf\[17\]\[12\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 rvsingle.dp.rf.rf\[19\]\[19\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 rvsingle.dp.rf.rf\[27\]\[17\] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 rvsingle.dp.rf.rf\[9\]\[18\] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 rvsingle.dp.rf.rf\[24\]\[12\] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 rvsingle.dp.rf.rf\[3\]\[21\] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold188 rvsingle.dp.rf.rf\[17\]\[18\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold199 rvsingle.dp.rf.rf\[19\]\[17\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _04738_ _04733_ _04725_ _04739_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _04628_ _04631_ _04675_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__a21oi_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ PC[22] _04597_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__nor2_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ _01469_ rvsingle.dp.rf.rf\[26\]\[22\] VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__or2_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _01248_ _03586_ _03597_ _03645_ _03647_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__a32o_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _01694_ _03574_ _03578_ _01221_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__o211ai_2
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _02504_ _01083_ _02505_ _02529_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__nand4_4
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _03507_ _01702_ _03509_ _01446_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_166_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10620_ _05209_ rvsingle.dp.rf.rf\[22\]\[13\] _05205_ VGND VGND VPWR VPWR _05210_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10551_ _05170_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10482_ _05128_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13270_ clknet_leaf_62_clk _00728_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12221_ _06068_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12152_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11103_ _05187_ net311 _05469_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__mux2_1
X_12083_ _05724_ net540 _06010_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__mux2_1
X_11034_ _05307_ net657 _05443_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__mux2_1
X_12985_ clknet_leaf_9_clk _00443_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11936_ _05932_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11867_ _05895_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10818_ _05322_ net638 _05320_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11798_ net32 VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10749_ _04774_ rvsingle.dp.rf.rf\[20\]\[7\] _05274_ VGND VGND VPWR VPWR _05281_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xload_slew1 DataAdr[16] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12419_ clknet_leaf_115_clk _00903_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13399_ clknet_leaf_6_clk _00827_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07960_ rvsingle.dp.rf.rf\[12\]\[0\] _01619_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_4_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_06911_ _01208_ _01825_ _01831_ _01478_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__o211ai_1
X_07891_ rvsingle.dp.rf.rf\[11\]\[2\] _01901_ _02811_ VGND VGND VPWR VPWR _02812_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09630_ PC[10] _04475_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__xor2_4
X_06842_ _01381_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__buf_8
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06773_ _01444_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__buf_6
X_09561_ _04414_ _04415_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__or2_1
X_08512_ _02117_ rvsingle.dp.rf.rf\[8\]\[13\] _03432_ _01542_ VGND VGND VPWR VPWR
+ _03433_ sky130_fd_sc_hd__o211ai_1
X_09492_ _02150_ VGND VGND VPWR VPWR WriteData[17] sky130_fd_sc_hd__inv_2
XFILLER_0_65_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08443_ _03352_ _03363_ _01682_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__nand3_2
XFILLER_0_148_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08374_ _03291_ _03292_ _01721_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07325_ rvsingle.dp.rf.rf\[15\]\[16\] _01509_ _01491_ VGND VGND VPWR VPWR _02246_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07256_ rvsingle.dp.rf.rf\[20\]\[17\] rvsingle.dp.rf.rf\[21\]\[17\] rvsingle.dp.rf.rf\[22\]\[17\]
+ rvsingle.dp.rf.rf\[23\]\[17\] _02176_ _01696_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06207_ _01130_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__buf_8
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07187_ _01666_ rvsingle.dp.rf.rf\[28\]\[17\] VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06138_ Instr[3] Instr[2] VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__nor2_4
XFILLER_0_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09828_ PC[24] PC[25] _04659_ PC[26] VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__a31o_1
X_09759_ PC[20] PC[21] _04582_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__and3_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ clknet_leaf_140_clk _00228_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _05820_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__clkbuf_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _05757_ net250 _05775_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10603_ _04770_ rvsingle.dp.rf.rf\[22\]\[6\] _05194_ VGND VGND VPWR VPWR _05200_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11583_ _05439_ net541 _05729_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13322_ clknet_leaf_104_clk _00780_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10534_ net78 _05155_ _05161_ _05157_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13253_ clknet_leaf_121_clk _00711_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10465_ net166 _05103_ _05119_ _04970_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12204_ _05898_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13184_ clknet_leaf_13_clk _00642_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10396_ _04814_ net480 _05071_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__mux2_1
X_12135_ _04876_ _04726_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12066_ _04876_ net466 _05994_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__mux2_1
X_11017_ _05295_ rvsingle.dp.rf.rf\[31\]\[19\] _05431_ VGND VGND VPWR VPWR _05441_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12968_ clknet_leaf_105_clk _00426_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11919_ _05923_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ clknet_leaf_116_clk _00357_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07110_ _01258_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__buf_6
XFILLER_0_126_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08090_ rvsingle.dp.rf.rf\[9\]\[1\] _01645_ _01667_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07041_ _01150_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__buf_12
XFILLER_0_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08992_ rvsingle.dp.rf.rf\[28\]\[27\] rvsingle.dp.rf.rf\[29\]\[27\] _01193_ VGND
+ VGND VPWR VPWR _03912_ sky130_fd_sc_hd__mux2_1
X_07943_ rvsingle.dp.rf.rf\[1\]\[0\] _01675_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07874_ _02792_ _02410_ _02794_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__nand3_1
X_09613_ Instr[27] PC[7] _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__a21oi_1
X_06825_ rvsingle.dp.rf.rf\[13\]\[23\] _01646_ _01520_ VGND VGND VPWR VPWR _01746_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_97_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09544_ _01114_ net825 _04397_ _02800_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06756_ _01645_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__buf_6
XFILLER_0_39_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09475_ _04378_ VGND VGND VPWR VPWR WriteData[0] sky130_fd_sc_hd__clkbuf_4
X_06687_ rvsingle.dp.rf.rf\[11\]\[20\] _01607_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08426_ _02005_ rvsingle.dp.rf.rf\[26\]\[9\] _01104_ VGND VGND VPWR VPWR _03347_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08357_ _01531_ _03274_ _03275_ _02410_ _03277_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07308_ rvsingle.dp.rf.rf\[29\]\[16\] _01540_ _01543_ VGND VGND VPWR VPWR _02229_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08288_ rvsingle.dp.rf.rf\[27\]\[10\] _01255_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07239_ rvsingle.dp.rf.rf\[12\]\[17\] rvsingle.dp.rf.rf\[13\]\[17\] rvsingle.dp.rf.rf\[14\]\[17\]
+ rvsingle.dp.rf.rf\[15\]\[17\] _01192_ _01728_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10250_ _04814_ net730 _04989_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10181_ _04853_ net464 _04952_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12822_ clknet_leaf_31_clk _00280_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12753_ clknet_leaf_49_clk _00211_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _05811_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12684_ clknet_leaf_54_clk _00142_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ net107 _05778_ _05742_ _05501_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11566_ _04785_ _05732_ _05733_ _05060_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13305_ clknet_leaf_19_clk _00763_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10517_ _05150_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__buf_8
X_11497_ _05700_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13236_ clknet_leaf_58_clk _00694_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10448_ _04770_ rvsingle.dp.rf.rf\[24\]\[6\] _05103_ VGND VGND VPWR VPWR _05109_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13167_ clknet_leaf_49_clk _00625_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10379_ _05064_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__buf_6
X_12118_ _05173_ net642 _06019_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__mux2_1
X_13098_ clknet_leaf_82_clk _00556_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_12049_ _05992_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06610_ _01530_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__buf_6
X_07590_ _01518_ rvsingle.dp.rf.rf\[22\]\[4\] VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06541_ _01190_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06472_ _01089_ rvsingle.dp.rf.rf\[3\]\[28\] _01261_ _01393_ VGND VGND VPWR VPWR
+ _01394_ sky130_fd_sc_hd__o211a_1
X_09260_ _01411_ _01412_ _04176_ _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_146_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08211_ rvsingle.dp.rf.rf\[28\]\[11\] rvsingle.dp.rf.rf\[29\]\[11\] rvsingle.dp.rf.rf\[30\]\[11\]
+ rvsingle.dp.rf.rf\[31\]\[11\] _01730_ _01808_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__mux4_1
X_09191_ _01085_ WriteData[31] _01180_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08142_ _02476_ _03058_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08073_ _02990_ _02991_ _02273_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07024_ rvsingle.dp.rf.rf\[11\]\[19\] _01943_ _01944_ VGND VGND VPWR VPWR _01945_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08975_ rvsingle.dp.rf.rf\[13\]\[25\] _01297_ _01310_ _03894_ VGND VGND VPWR VPWR
+ _03895_ sky130_fd_sc_hd__o211ai_1
Xhold15 rvsingle.dp.rf.rf\[0\]\[10\] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 rvsingle.dp.rf.rf\[27\]\[20\] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 rvsingle.dp.rf.rf\[7\]\[3\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _02831_ _02836_ _01187_ _02846_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__o211ai_4
Xhold48 rvsingle.dp.rf.rf\[10\]\[31\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 rvsingle.dp.rf.rf\[13\]\[31\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ rvsingle.dp.rf.rf\[29\]\[2\] _01508_ _02395_ _02777_ VGND VGND VPWR VPWR
+ _02778_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06808_ rvsingle.dp.rf.rf\[24\]\[20\] rvsingle.dp.rf.rf\[25\]\[20\] rvsingle.dp.rf.rf\[26\]\[20\]
+ rvsingle.dp.rf.rf\[27\]\[20\] _01726_ _01728_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07788_ _02703_ _02491_ _02708_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__nand3_1
X_09527_ _04121_ _04122_ _03731_ _04211_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__or4_4
XFILLER_0_149_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06739_ _01604_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09458_ _04364_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__buf_6
XFILLER_0_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08409_ _01268_ rvsingle.dp.rf.rf\[0\]\[9\] VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09389_ _04165_ _04237_ _03774_ _03831_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11420_ _05207_ net367 _05657_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11351_ _05209_ rvsingle.dp.rf.rf\[14\]\[13\] _05618_ VGND VGND VPWR VPWR _05621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10302_ _05027_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11282_ _05583_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13021_ clknet_leaf_145_clk _00479_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10233_ _04977_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__buf_6
X_10164_ _04808_ net415 _04941_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__mux2_1
X_10095_ _04893_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12805_ clknet_leaf_123_clk _00263_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10997_ _05385_ net455 _05419_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12736_ clknet_leaf_116_clk _00194_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12667_ clknet_leaf_141_clk _00125_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11618_ _04973_ _05457_ net109 VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12598_ clknet_leaf_33_clk _00056_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11549_ _04967_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold507 rvsingle.dp.rf.rf\[22\]\[19\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold518 rvsingle.dp.rf.rf\[19\]\[30\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 rvsingle.dp.rf.rf\[18\]\[4\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13219_ clknet_leaf_125_clk _00677_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _01498_ rvsingle.dp.rf.rf\[12\]\[15\] VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__or2_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ _02622_ _02625_ _02364_ _02631_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_73_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08691_ _01567_ rvsingle.dp.rf.rf\[18\]\[14\] _02031_ _03611_ VGND VGND VPWR VPWR
+ _03612_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_73_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07642_ _02163_ rvsingle.dp.rf.rf\[20\]\[4\] VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07573_ rvsingle.dp.rf.rf\[11\]\[4\] _02478_ _01523_ VGND VGND VPWR VPWR _02494_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09312_ _04225_ _04136_ _04227_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__nand3_4
XFILLER_0_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06524_ _01444_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09243_ _03572_ _03755_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06455_ _01376_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09174_ rvsingle.dp.rf.rf\[20\]\[31\] rvsingle.dp.rf.rf\[21\]\[31\] rvsingle.dp.rf.rf\[22\]\[31\]
+ rvsingle.dp.rf.rf\[23\]\[31\] _02212_ _01120_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__mux4_1
X_06386_ _01307_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08125_ net822 _03045_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__nand2_2
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ rvsingle.dp.rf.rf\[5\]\[1\] _02271_ _01436_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07007_ _01581_ _01897_ _01837_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08958_ _02212_ _01962_ _03855_ _03878_ VGND VGND VPWR VPWR WriteData[25] sky130_fd_sc_hd__o211a_4
X_07909_ rvsingle.dp.rf.rf\[21\]\[2\] _02275_ _01436_ _02829_ VGND VGND VPWR VPWR
+ _02830_ sky130_fd_sc_hd__o211ai_1
X_08889_ rvsingle.dp.rf.rf\[28\]\[24\] rvsingle.dp.rf.rf\[29\]\[24\] rvsingle.dp.rf.rf\[30\]\[24\]
+ rvsingle.dp.rf.rf\[31\]\[24\] _01463_ _01471_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10920_ _04785_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__clkbuf_4
X_10851_ _04814_ _05316_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__nand2_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10782_ _05299_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__clkbuf_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ clknet_leaf_96_clk _01005_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12452_ clknet_leaf_107_clk _00936_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11403_ _05377_ rvsingle.dp.rf.rf\[13\]\[4\] _05646_ VGND VGND VPWR VPWR _05650_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12383_ clknet_leaf_132_clk _00867_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11334_ _05534_ rvsingle.dp.rf.rf\[14\]\[5\] _05607_ VGND VGND VPWR VPWR _05612_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11265_ _05574_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13004_ clknet_leaf_51_clk _00462_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10216_ _04977_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__buf_8
X_11196_ _05536_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__clkbuf_1
X_10147_ _04770_ net656 _04930_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10078_ _04878_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12719_ clknet_leaf_27_clk _00177_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06240_ _01161_ _01094_ _01134_ _01163_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_128_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06171_ Instr[20] VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold304 rvsingle.dp.rf.rf\[2\]\[22\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 rvsingle.dp.rf.rf\[26\]\[10\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 rvsingle.dp.rf.rf\[21\]\[30\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold337 rvsingle.dp.rf.rf\[26\]\[30\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 rvsingle.dp.rf.rf\[0\]\[24\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09930_ _04426_ _04406_ _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_22_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold359 rvsingle.dp.rf.rf\[7\]\[29\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _04398_ _04683_ _04690_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[29\] sky130_fd_sc_hd__o21ai_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _01202_ _01351_ _03713_ _03726_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__o211ai_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _04585_ _04625_ _04609_ _04626_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__or4_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ rvsingle.dp.rf.rf\[29\]\[15\] _02627_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _03592_ _01716_ _01460_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__a211o_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _01690_ rvsingle.dp.rf.rf\[0\]\[4\] VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__or2_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_867 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07556_ _01518_ rvsingle.dp.rf.rf\[2\]\[4\] VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06507_ _01426_ rvsingle.dp.rf.rf\[30\]\[21\] _01427_ VGND VGND VPWR VPWR _01428_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07487_ _01545_ rvsingle.dp.rf.rf\[12\]\[6\] VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09226_ _01480_ _01453_ _01582_ _01579_ _01739_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__o41a_1
XFILLER_0_63_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06438_ _01232_ _01355_ _01359_ _01224_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09157_ rvsingle.dp.rf.rf\[16\]\[31\] rvsingle.dp.rf.rf\[17\]\[31\] rvsingle.dp.rf.rf\[18\]\[31\]
+ rvsingle.dp.rf.rf\[19\]\[31\] _01225_ _01226_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__mux4_1
X_06369_ rvsingle.dp.rf.rf\[4\]\[29\] rvsingle.dp.rf.rf\[5\]\[29\] rvsingle.dp.rf.rf\[6\]\[29\]
+ rvsingle.dp.rf.rf\[7\]\[29\] _01195_ _01202_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__mux4_1
X_08108_ _01880_ _03025_ _03026_ _01599_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09088_ _01209_ _04003_ _01223_ _04007_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_20_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08039_ _02952_ _02954_ _01216_ _02959_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__o211ai_1
X_11050_ _05459_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__buf_6
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10001_ _04505_ _04506_ _04544_ _04812_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__a31o_4
X_11952_ _05942_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10903_ _05375_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__clkbuf_1
X_11883_ _05531_ rvsingle.dp.rf.rf\[6\]\[3\] _05902_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10834_ _04781_ _04726_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10765_ _05289_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12504_ clknet_leaf_34_clk _00988_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10696_ _05251_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12435_ clknet_leaf_33_clk _00919_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12366_ clknet_leaf_71_clk _00850_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11317_ _05601_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__clkbuf_1
X_12297_ _06098_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__buf_6
X_11248_ _05364_ _05365_ _05525_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__o21ai_1
X_11179_ _04925_ _05061_ net74 VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07410_ _02117_ rvsingle.dp.rf.rf\[10\]\[7\] _01654_ _02330_ VGND VGND VPWR VPWR
+ _02331_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08390_ _01188_ _03297_ _03310_ _01247_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__o211a_2
XFILLER_0_169_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07341_ _02256_ _01084_ _01153_ _02234_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__nand4_2
XFILLER_0_58_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07272_ rvsingle.dp.rf.rf\[26\]\[16\] rvsingle.dp.rf.rf\[27\]\[16\] _01726_ VGND
+ VGND VPWR VPWR _02193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09011_ rvsingle.dp.rf.rf\[4\]\[27\] rvsingle.dp.rf.rf\[5\]\[27\] rvsingle.dp.rf.rf\[6\]\[27\]
+ rvsingle.dp.rf.rf\[7\]\[27\] _01336_ _01451_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06223_ _01146_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__buf_8
XFILLER_0_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06154_ _01077_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__buf_4
Xhold101 rvsingle.dp.rf.rf\[7\]\[11\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold112 rvsingle.dp.rf.rf\[31\]\[0\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 rvsingle.dp.rf.rf\[16\]\[9\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold134 rvsingle.dp.rf.rf\[5\]\[26\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold145 rvsingle.dp.rf.rf\[1\]\[21\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 rvsingle.dp.rf.rf\[27\]\[19\] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 rvsingle.dp.rf.rf\[17\]\[10\] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ Instr[8] VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__clkbuf_2
Xhold178 rvsingle.dp.rf.rf\[13\]\[0\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 rvsingle.dp.rf.rf\[19\]\[11\] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _04644_ _04653_ _04667_ _04634_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__or4_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _04611_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__buf_2
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06987_ rvsingle.dp.rf.rf\[28\]\[22\] rvsingle.dp.rf.rf\[29\]\[22\] rvsingle.dp.rf.rf\[30\]\[22\]
+ rvsingle.dp.rf.rf\[31\]\[22\] _01329_ _01456_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__mux4_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _03646_ _01183_ _02261_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__nand3_2
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _03575_ _01716_ _01460_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07608_ _02516_ _01146_ _02528_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__nand3_4
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08588_ rvsingle.dp.rf.rf\[23\]\[12\] _01901_ _03508_ VGND VGND VPWR VPWR _03509_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07539_ _02456_ _02457_ _01444_ _02459_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10550_ _04814_ net372 _05151_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09209_ _01060_ _04120_ _04123_ _04124_ _04127_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__o32a_1
X_10481_ _04840_ net626 _05126_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12220_ _06068_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12151_ _04722_ _04723_ _04724_ _05003_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__or4_1
X_11102_ _04898_ _05183_ _05457_ _05483_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12082_ _06009_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__buf_6
Xhold690 rvsingle.dp.rf.rf\[11\]\[16\] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__dlygate4sd3_1
X_11033_ _05449_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12984_ clknet_leaf_23_clk _00442_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11935_ _05763_ net292 _05924_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__mux2_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _05639_ net266 _05885_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__mux2_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10817_ _04746_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__buf_2
XFILLER_0_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11797_ _05857_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10748_ _05280_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10679_ _05242_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12418_ clknet_leaf_130_clk _00902_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_13398_ clknet_leaf_31_clk _00826_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12349_ _06126_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06910_ _01826_ _01309_ _01229_ _01830_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__a211o_1
X_07890_ _01903_ rvsingle.dp.rf.rf\[10\]\[2\] _01243_ VGND VGND VPWR VPWR _02811_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06841_ _01619_ rvsingle.dp.rf.rf\[4\]\[23\] _01654_ VGND VGND VPWR VPWR _01762_
+ sky130_fd_sc_hd__o21bai_1
X_09560_ PC[4] _02532_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__nor2_1
X_06772_ rvsingle.dp.rf.rf\[13\]\[20\] _01688_ _01689_ _01692_ VGND VGND VPWR VPWR
+ _01693_ sky130_fd_sc_hd__o211ai_1
X_08511_ rvsingle.dp.rf.rf\[9\]\[13\] _01096_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__or2b_1
X_09491_ _02065_ VGND VGND VPWR VPWR WriteData[18] sky130_fd_sc_hd__inv_6
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08442_ _03355_ _03357_ _01853_ _03362_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08373_ rvsingle.dp.rf.rf\[11\]\[8\] _01424_ _03293_ VGND VGND VPWR VPWR _03294_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07324_ _01269_ rvsingle.dp.rf.rf\[14\]\[16\] VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07255_ _01425_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__buf_8
XFILLER_0_116_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06206_ Instr[22] VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__inv_2
X_07186_ _02103_ _02104_ _02106_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06137_ Instr[6] Instr[4] VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09827_ PC[24] PC[25] PC[26] _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__and4_1
X_09758_ _04594_ _04452_ _04596_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[20\] sky130_fd_sc_hd__o21ai_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08709_ _03627_ _02488_ _03629_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__nand3_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ PC[14] _04522_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__xor2_2
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _05757_ net584 _05817_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11651_ net200 _05778_ _05756_ _05457_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10602_ _05199_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11582_ net163 _05726_ _05751_ _05737_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13321_ clknet_leaf_99_clk _00779_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10533_ _05113_ _05114_ _05115_ _05061_ _04773_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__o311a_1
XFILLER_0_135_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13252_ clknet_leaf_19_clk _00710_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10464_ _05113_ _05114_ _05115_ _04924_ _04795_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__o311a_1
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ _05898_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13183_ clknet_leaf_144_clk _00641_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10395_ _05079_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12134_ _06037_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12065_ _06000_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11016_ _05440_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ clknet_leaf_98_clk _00425_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _04839_ net665 _05913_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12898_ clknet_leaf_141_clk _00356_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ _05886_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_998 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07040_ net822 VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__buf_8
XFILLER_0_42_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08991_ rvsingle.dp.rf.rf\[24\]\[27\] rvsingle.dp.rf.rf\[25\]\[27\] rvsingle.dp.rf.rf\[26\]\[27\]
+ rvsingle.dp.rf.rf\[27\]\[27\] _01330_ _01302_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07942_ rvsingle.dp.rf.rf\[0\]\[0\] _01256_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07873_ _01558_ rvsingle.dp.rf.rf\[22\]\[2\] _01259_ _02793_ VGND VGND VPWR VPWR
+ _02794_ sky130_fd_sc_hd__o211ai_1
X_09612_ _04448_ PC[6] Instr[26] VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__and3_1
X_06824_ _01744_ rvsingle.dp.rf.rf\[12\]\[23\] VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09543_ _04371_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__nand2_1
X_06755_ rvsingle.dp.rf.rf\[19\]\[20\] _01675_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__and2b_1
XFILLER_0_148_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09474_ _04377_ _02885_ _02906_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__and3_2
XFILLER_0_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06686_ _01606_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__buf_6
X_08425_ _03342_ _03343_ _03345_ _01632_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_149_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08356_ _01545_ rvsingle.dp.rf.rf\[22\]\[8\] _02031_ _03276_ VGND VGND VPWR VPWR
+ _03277_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07307_ _01383_ rvsingle.dp.rf.rf\[28\]\[16\] VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__nor2_1
X_08287_ _03206_ _03207_ _02483_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07238_ _02156_ _01717_ _01461_ _02158_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07169_ rvsingle.dp.rf.rf\[25\]\[18\] _01943_ _01717_ _02089_ VGND VGND VPWR VPWR
+ _02090_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_14_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10180_ _04953_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12821_ clknet_leaf_26_clk _00279_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12752_ clknet_leaf_52_clk _00210_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11703_ _04813_ net552 _05806_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ clknet_leaf_88_clk _00141_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11634_ _05780_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11565_ net14 _05726_ _05742_ _05737_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13304_ clknet_leaf_26_clk _00762_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10516_ Instr[8] _04732_ _05149_ Instr[7] VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__or4b_1
XFILLER_0_123_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11496_ _04813_ net338 _05695_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13235_ clknet_leaf_47_clk _00693_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10447_ _05108_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13166_ clknet_leaf_53_clk _00624_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10378_ _04988_ _05068_ _05069_ _05065_ net75 VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12117_ _06028_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13097_ clknet_leaf_92_clk _00555_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_12048_ _04823_ net357 _05983_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06540_ _01460_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__buf_6
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06471_ _01099_ rvsingle.dp.rf.rf\[2\]\[28\] VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_190 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08210_ _03126_ _03129_ _03130_ _01694_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__o22ai_2
X_09190_ _01378_ _04093_ _04099_ _04109_ _01154_ VGND VGND VPWR VPWR WriteData[31]
+ sky130_fd_sc_hd__o311a_4
XFILLER_0_90_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08141_ _02377_ _02374_ _02464_ _03061_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08072_ rvsingle.dp.rf.rf\[29\]\[1\] _02275_ _01436_ _02992_ VGND VGND VPWR VPWR
+ _02993_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07023_ _01242_ rvsingle.dp.rf.rf\[10\]\[19\] _01728_ VGND VGND VPWR VPWR _01944_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08974_ _01193_ rvsingle.dp.rf.rf\[12\]\[25\] VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__or2_1
Xhold16 rvsingle.dp.rf.rf\[16\]\[20\] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 rvsingle.dp.rf.rf\[9\]\[22\] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _01702_ _02838_ _02840_ _02845_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__o31ai_2
Xhold38 rvsingle.dp.rf.rf\[12\]\[31\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 rvsingle.dp.rf.rf\[8\]\[31\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07856_ _01877_ rvsingle.dp.rf.rf\[28\]\[2\] VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__or2_1
X_06807_ _01727_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__clkbuf_8
X_07787_ _02704_ _02705_ _02706_ _02707_ _01111_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__o221ai_2
X_09526_ _04273_ VGND VGND VPWR VPWR DataAdr[14] sky130_fd_sc_hd__inv_6
X_06738_ rvsingle.dp.rf.rf\[25\]\[20\] _01658_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09457_ _04140_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__buf_4
XFILLER_0_164_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06669_ _01583_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__nand2_1
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08408_ _03321_ _03323_ _02527_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_19_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09388_ _03775_ _03831_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08339_ rvsingle.dp.rf.rf\[31\]\[8\] _01677_ _03259_ VGND VGND VPWR VPWR _03260_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11350_ _05620_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10301_ _04765_ net545 _05022_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11281_ _05209_ rvsingle.dp.rf.rf\[15\]\[13\] _05580_ VGND VGND VPWR VPWR _05583_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13020_ clknet_leaf_13_clk _00478_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10232_ net106 _04978_ _04988_ _04985_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__a22o_1
X_10163_ _04944_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
X_10094_ _04892_ net228 _04847_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12804_ clknet_leaf_123_clk _00262_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10996_ _05429_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ clknet_leaf_2_clk _00193_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12666_ clknet_leaf_3_clk _00124_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11617_ _04720_ _05367_ _04967_ _04968_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__and4_2
XFILLER_0_5_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12597_ clknet_leaf_37_clk _00055_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11548_ _04968_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold508 rvsingle.dp.rf.rf\[15\]\[26\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 rvsingle.dp.rf.rf\[2\]\[12\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11479_ _05381_ rvsingle.dp.rf.rf\[12\]\[7\] _05684_ VGND VGND VPWR VPWR _05691_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13218_ clknet_leaf_137_clk _00676_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ clknet_leaf_143_clk _00607_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _01520_ _02626_ _02628_ _01564_ _02630_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__o311ai_2
X_08690_ rvsingle.dp.rf.rf\[19\]\[14\] _01779_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__or2b_1
X_07641_ rvsingle.dp.rf.rf\[16\]\[4\] rvsingle.dp.rf.rf\[17\]\[4\] rvsingle.dp.rf.rf\[18\]\[4\]
+ rvsingle.dp.rf.rf\[19\]\[4\] _02176_ _02162_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__mux4_1
X_07572_ _01493_ rvsingle.dp.rf.rf\[10\]\[4\] VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09311_ _04220_ _04223_ _04226_ _03650_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06523_ _01172_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__buf_8
XFILLER_0_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09242_ _03231_ _04160_ _03753_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06454_ _01145_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09173_ _01114_ _04088_ _01118_ _04092_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__o211a_1
X_06385_ _01306_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08124_ _01856_ net825 _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_114_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08055_ _01695_ rvsingle.dp.rf.rf\[4\]\[1\] VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07006_ _01898_ _01925_ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08957_ _03861_ _03866_ _01378_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_76_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07908_ _01349_ rvsingle.dp.rf.rf\[20\]\[2\] VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__or2_1
X_08888_ _03805_ _03807_ _01722_ _03808_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__o2bb2a_1
X_07839_ rvsingle.dp.rf.rf\[15\]\[2\] _01539_ _02759_ VGND VGND VPWR VPWR _02760_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10850_ _05085_ _05342_ _05325_ net98 VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09509_ _02662_ VGND VGND VPWR VPWR WriteData[5] sky130_fd_sc_hd__inv_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10781_ _04846_ net571 _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__mux2_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12520_ clknet_leaf_106_clk _01004_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ clknet_leaf_126_clk _00935_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11402_ _05649_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12382_ clknet_leaf_133_clk _00866_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_90 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11333_ _05611_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11264_ _05534_ net741 _05569_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13003_ clknet_leaf_89_clk _00461_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10215_ _04724_ _04927_ _04975_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__or4_4
X_11195_ _05496_ net757 _05528_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__mux2_1
X_10146_ _04935_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10077_ _04877_ net223 _04847_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10979_ _05420_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12718_ clknet_leaf_71_clk _00176_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12649_ clknet_leaf_95_clk _00107_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06170_ _01093_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__buf_4
XFILLER_0_170_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold305 rvsingle.dp.rf.rf\[30\]\[27\] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 rvsingle.dp.rf.rf\[5\]\[20\] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold327 rvsingle.dp.rf.rf\[4\]\[18\] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold338 rvsingle.dp.rf.rf\[12\]\[15\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 rvsingle.dp.rf.rf\[18\]\[17\] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09860_ _04366_ _04688_ _04689_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__nand3_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _01587_ _03730_ _01486_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__a21oi_1
X_09791_ _04619_ _04620_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__nand2_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ rvsingle.dp.rf.rf\[31\]\[15\] _01487_ _01523_ VGND VGND VPWR VPWR _03663_
+ sky130_fd_sc_hd__o21ai_1
X_08673_ _02450_ rvsingle.dp.rf.rf\[30\]\[14\] _01427_ _03593_ VGND VGND VPWR VPWR
+ _03594_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07624_ rvsingle.dp.rf.rf\[3\]\[4\] _02288_ _02544_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ _02374_ _02377_ _02464_ _02468_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_49_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06506_ _01197_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07486_ _02405_ _02406_ _01131_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09225_ _01834_ _01838_ _04143_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__o21ai_2
X_06437_ _01356_ _01311_ _01209_ _01358_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09156_ _01189_ _04069_ _04075_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06368_ _01289_ _01184_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__nand2_2
XFILLER_0_161_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08107_ _01769_ rvsingle.dp.rf.rf\[18\]\[1\] _01604_ _03027_ VGND VGND VPWR VPWR
+ _03028_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_16_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09087_ _01201_ _04004_ _04006_ _01915_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_110_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_110_clk sky130_fd_sc_hd__clkbuf_16
X_06299_ _01221_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__buf_6
XFILLER_0_102_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08038_ _02955_ _02956_ _01172_ _02958_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10000_ _01169_ _02259_ _01170_ _04810_ _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__o32a_1
XFILLER_0_101_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09989_ _04802_ net648 _04791_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11951_ _05728_ rvsingle.dp.rf.rf\[4\]\[2\] _05940_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__mux2_1
X_10902_ _05322_ rvsingle.dp.rf.rf\[18\]\[2\] _05373_ VGND VGND VPWR VPWR _05375_
+ sky130_fd_sc_hd__mux2_1
X_11882_ _05904_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10833_ _05331_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10764_ _04808_ net647 _05285_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12503_ clknet_leaf_6_clk _00987_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10695_ _05212_ net500 _05246_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12434_ clknet_leaf_36_clk _00918_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12365_ clknet_leaf_44_clk _00849_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_101_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_101_clk sky130_fd_sc_hd__clkbuf_16
X_11316_ _05187_ net407 _05591_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12296_ _04728_ _04925_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__nand2_2
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11247_ net80 VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__inv_2
X_11178_ _04916_ _04918_ _04922_ _05058_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__and4_2
X_10129_ _04920_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__buf_4
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07340_ _01483_ net824 _01177_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07271_ rvsingle.dp.rf.rf\[28\]\[16\] rvsingle.dp.rf.rf\[29\]\[16\] rvsingle.dp.rf.rf\[30\]\[16\]
+ rvsingle.dp.rf.rf\[31\]\[16\] _01242_ _01434_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09010_ _03926_ _03928_ _02191_ _03929_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_73_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06222_ _01145_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06153_ _01076_ _01071_ _01062_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__nand3_1
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold102 rvsingle.dp.rf.rf\[11\]\[24\] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold113 rvsingle.dp.rf.rf\[11\]\[4\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 rvsingle.dp.rf.rf\[14\]\[0\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold135 rvsingle.dp.rf.rf\[17\]\[7\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold146 rvsingle.dp.rf.rf\[25\]\[19\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 rvsingle.dp.rf.rf\[11\]\[13\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold168 rvsingle.dp.rf.rf\[8\]\[12\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold179 rvsingle.dp.rf.rf\[17\]\[26\] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _04737_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__clkbuf_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ PC[24] PC[25] PC[26] PC[27] _04617_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__o41a_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06986_ _01208_ _01899_ _01906_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__o21bai_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ PC[20] PC[21] PC[22] _04582_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__and4_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _02505_ _03643_ _03620_ _02375_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__a31o_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _01423_ rvsingle.dp.rf.rf\[15\]\[14\] _01427_ _03576_ VGND VGND VPWR VPWR
+ _03577_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07607_ _02521_ _02526_ _02527_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__nand3_1
XFILLER_0_135_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _01903_ rvsingle.dp.rf.rf\[22\]\[12\] _01243_ VGND VGND VPWR VPWR _03508_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07538_ rvsingle.dp.rf.rf\[23\]\[6\] _02288_ _02458_ VGND VGND VPWR VPWR _02459_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07469_ _01847_ rvsingle.dp.rf.rf\[16\]\[6\] VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09208_ _04121_ _04122_ _01066_ _04125_ _04126_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__o32a_1
XFILLER_0_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10480_ _05127_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09139_ _03775_ _03910_ _04056_ _04058_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_122_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12150_ _05721_ _06045_ _06046_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11101_ _05084_ _05371_ net652 VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__o21a_1
X_12081_ _04737_ _04919_ _04733_ _04725_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__or4b_2
Xhold680 rvsingle.dp.rf.rf\[4\]\[12\] VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold691 rvsingle.dp.rf.rf\[23\]\[26\] VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ _05407_ net502 _05443_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12983_ clknet_leaf_9_clk _00441_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11934_ _05931_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _05894_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__clkbuf_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10816_ _05321_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11796_ _05639_ net699 _05836_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10747_ _04770_ rvsingle.dp.rf.rf\[20\]\[6\] _05274_ VGND VGND VPWR VPWR _05280_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10678_ _04774_ net318 _05235_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12417_ clknet_leaf_140_clk _00901_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13397_ clknet_leaf_37_clk _00825_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12348_ _04869_ net475 _06121_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12279_ _04869_ net620 _06073_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06840_ _01758_ _01559_ _01759_ _01760_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__a211oi_1
X_06771_ _01691_ rvsingle.dp.rf.rf\[12\]\[20\] VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08510_ rvsingle.dp.rf.rf\[11\]\[13\] _01860_ _01259_ VGND VGND VPWR VPWR _03431_
+ sky130_fd_sc_hd__o21ai_1
X_09490_ _02011_ VGND VGND VPWR VPWR WriteData[19] sky130_fd_sc_hd__inv_2
XFILLER_0_77_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08441_ _01605_ _03358_ _03359_ _01511_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08372_ _01426_ rvsingle.dp.rf.rf\[10\]\[8\] _01427_ VGND VGND VPWR VPWR _03293_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07323_ _01132_ _02241_ _02243_ _01526_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07254_ rvsingle.dp.rf.rf\[16\]\[17\] rvsingle.dp.rf.rf\[17\]\[17\] rvsingle.dp.rf.rf\[18\]\[17\]
+ rvsingle.dp.rf.rf\[19\]\[17\] _01329_ _01456_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06205_ rvsingle.dp.rf.rf\[12\]\[30\] rvsingle.dp.rf.rf\[13\]\[30\] _01128_ VGND
+ VGND VPWR VPWR _01129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07185_ _01848_ rvsingle.dp.rf.rf\[24\]\[17\] _02105_ _01759_ VGND VGND VPWR VPWR
+ _02106_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_42_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06136_ Instr[12] Instr[13] VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09826_ PC[22] PC[23] _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__and3_1
X_09757_ _04422_ _04423_ _04595_ _04427_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__o211ai_1
X_06969_ _01098_ rvsingle.dp.rf.rf\[22\]\[22\] VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__nor2_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08708_ rvsingle.dp.rf.rf\[15\]\[14\] _02481_ _03628_ VGND VGND VPWR VPWR _03629_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09688_ _04531_ _04532_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__or2_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _03548_ _01146_ _03559_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__nand3_4
XFILLER_0_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _05783_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__clkbuf_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10601_ _04765_ rvsingle.dp.rf.rf\[22\]\[5\] _05194_ VGND VGND VPWR VPWR _05199_
+ sky130_fd_sc_hd__mux2_1
X_11581_ _04823_ _05732_ _05733_ _05097_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10532_ _05160_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__clkbuf_1
X_13320_ clknet_leaf_121_clk _00778_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13251_ clknet_leaf_130_clk _00709_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10463_ _05118_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12202_ _06066_ _06045_ _06067_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__o21ai_1
X_13182_ clknet_leaf_147_clk _00640_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10394_ _04808_ net523 _05071_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__mux2_1
X_12133_ _04869_ net482 _06031_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12064_ _04869_ net727 _05994_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11015_ _05439_ rvsingle.dp.rf.rf\[31\]\[18\] _05431_ VGND VGND VPWR VPWR _05440_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12966_ clknet_leaf_114_clk _00424_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _05922_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__clkbuf_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ clknet_leaf_140_clk _00355_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _04845_ net811 _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11779_ _05849_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08990_ _03831_ _03908_ _03909_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__and3_2
X_07941_ _02851_ _02803_ _02856_ _02751_ _02861_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__o2111a_1
X_07872_ rvsingle.dp.rf.rf\[23\]\[2\] _01544_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__or2b_1
X_09611_ Instr[25] _04429_ _04439_ _04419_ _04461_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__o221ai_2
X_06823_ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__buf_8
X_09542_ _04368_ PC[0] _04369_ _04372_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__nand4_1
X_06754_ _01096_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06685_ Instr[20] VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09473_ _01154_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_90_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
X_08424_ _01562_ rvsingle.dp.rf.rf\[28\]\[9\] _03344_ _02485_ VGND VGND VPWR VPWR
+ _03345_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_164_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08355_ rvsingle.dp.rf.rf\[23\]\[8\] _01877_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07306_ _01383_ rvsingle.dp.rf.rf\[24\]\[16\] _02226_ _01543_ VGND VGND VPWR VPWR
+ _02227_ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08286_ rvsingle.dp.rf.rf\[25\]\[10\] _01797_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07237_ _01688_ rvsingle.dp.rf.rf\[7\]\[17\] _01456_ _02157_ VGND VGND VPWR VPWR
+ _02158_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07168_ _01417_ rvsingle.dp.rf.rf\[24\]\[18\] VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__or2_1
X_07099_ rvsingle.dp.rf.rf\[27\]\[18\] _01540_ _02019_ VGND VGND VPWR VPWR _02020_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09809_ PC[25] _04639_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12820_ clknet_leaf_64_clk _00278_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ clknet_leaf_37_clk _00209_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _05810_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ clknet_leaf_82_clk _00140_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _05740_ net332 _05775_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11564_ _04781_ _05732_ _05733_ _05097_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13303_ clknet_leaf_60_clk _00761_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10515_ _05148_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11495_ _05699_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10446_ _04765_ net765 _05103_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13234_ clknet_leaf_55_clk _00692_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10377_ _04987_ _05068_ _05069_ _05065_ net2 VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__a32o_1
X_13165_ clknet_leaf_90_clk _00623_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12116_ _04823_ net265 _06019_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__mux2_1
X_13096_ clknet_leaf_102_clk _00554_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12047_ _05991_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ clknet_leaf_36_clk _00407_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06470_ rvsingle.dp.rf.rf\[4\]\[28\] rvsingle.dp.rf.rf\[5\]\[28\] rvsingle.dp.rf.rf\[6\]\[28\]
+ rvsingle.dp.rf.rf\[7\]\[28\] _01099_ _01261_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_191 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08140_ _03060_ _02373_ _02317_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08071_ _01349_ rvsingle.dp.rf.rf\[28\]\[1\] VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07022_ _01424_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08973_ rvsingle.dp.rf.rf\[8\]\[25\] rvsingle.dp.rf.rf\[9\]\[25\] rvsingle.dp.rf.rf\[10\]\[25\]
+ rvsingle.dp.rf.rf\[11\]\[25\] _01330_ _01302_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 rvsingle.dp.rf.rf\[24\]\[0\] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 rvsingle.dp.rf.rf\[3\]\[0\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _02842_ _02844_ _01444_ _01216_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__a31oi_1
Xhold39 rvsingle.dp.rf.rf\[1\]\[17\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07855_ rvsingle.dp.rf.rf\[31\]\[2\] _01539_ _01520_ VGND VGND VPWR VPWR _02776_
+ sky130_fd_sc_hd__o21ai_1
X_06806_ _01197_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07786_ rvsingle.dp.rf.rf\[13\]\[3\] _01645_ _01667_ VGND VGND VPWR VPWR _02707_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09525_ _04268_ VGND VGND VPWR VPWR DataAdr[13] sky130_fd_sc_hd__inv_2
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06737_ _01557_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__buf_6
XFILLER_0_94_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06668_ _01179_ _01585_ _01586_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__o211ai_2
X_09456_ _04175_ _04190_ _04236_ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__nand4_4
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08407_ _01105_ _03324_ _03325_ _01511_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_149_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09387_ _03140_ net821 _04143_ _03112_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__o211ai_4
X_06599_ _01519_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__buf_8
XFILLER_0_35_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08338_ _03258_ rvsingle.dp.rf.rf\[30\]\[8\] _01604_ VGND VGND VPWR VPWR _03259_
+ sky130_fd_sc_hd__o21a_1
X_08269_ _01618_ rvsingle.dp.rf.rf\[6\]\[10\] _01551_ VGND VGND VPWR VPWR _03190_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10300_ _05026_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11280_ _05582_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10231_ _04981_ _04769_ _04982_ _04983_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__and4b_2
XFILLER_0_120_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10162_ _04802_ net504 _04941_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__mux2_1
X_10093_ _04891_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12803_ clknet_leaf_115_clk _00261_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_54_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10995_ _05428_ net644 _05419_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12734_ clknet_leaf_150_clk _00192_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12665_ clknet_leaf_8_clk _00123_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11616_ _05768_ _05722_ _05771_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12596_ clknet_leaf_58_clk _00054_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11547_ _05726_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__buf_6
XFILLER_0_80_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold509 rvsingle.dp.rf.rf\[13\]\[6\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11478_ _05690_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13217_ clknet_leaf_128_clk _00675_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10429_ _05095_ _05059_ _05096_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ clknet_leaf_147_clk _00606_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ clknet_leaf_10_clk _00537_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07640_ _02555_ _02560_ _01315_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07571_ _02487_ _02488_ _02490_ _02491_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_45_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
X_06522_ _01441_ rvsingle.dp.rf.rf\[23\]\[21\] _01301_ _01442_ VGND VGND VPWR VPWR
+ _01443_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09310_ _03729_ _03734_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06453_ _01351_ _01226_ _01361_ _01374_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__o211ai_2
X_09241_ _03313_ _03405_ _03748_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09172_ _01120_ _04089_ _01134_ _04091_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a211o_1
X_06384_ Instr[16] VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08123_ Instr[8] _01076_ _01071_ _01062_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__nand4_2
XFILLER_0_160_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08054_ rvsingle.dp.rf.rf\[0\]\[1\] rvsingle.dp.rf.rf\[1\]\[1\] rvsingle.dp.rf.rf\[2\]\[1\]
+ rvsingle.dp.rf.rf\[3\]\[1\] _02440_ _01470_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07005_ _01587_ _01897_ _01066_ _01075_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08956_ _01113_ _03871_ _03876_ _01117_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07907_ rvsingle.dp.rf.rf\[23\]\[2\] _01295_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__nor2_1
X_08887_ rvsingle.dp.rf.rf\[20\]\[24\] rvsingle.dp.rf.rf\[21\]\[24\] rvsingle.dp.rf.rf\[22\]\[24\]
+ rvsingle.dp.rf.rf\[23\]\[24\] _01469_ _01728_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07838_ _02627_ rvsingle.dp.rf.rf\[14\]\[2\] _01519_ VGND VGND VPWR VPWR _02759_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1000 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07769_ rvsingle.dp.rf.rf\[28\]\[3\] rvsingle.dp.rf.rf\[29\]\[3\] _01419_ VGND VGND
+ VPWR VPWR _02690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
X_09508_ _02427_ VGND VGND VPWR VPWR WriteData[6] sky130_fd_sc_hd__inv_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10780_ _05273_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__buf_8
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ _04153_ _02577_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand2_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12450_ clknet_leaf_128_clk _00934_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11401_ _05531_ rvsingle.dp.rf.rf\[13\]\[3\] _05646_ VGND VGND VPWR VPWR _05649_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12381_ clknet_leaf_135_clk _00865_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_80 ReadData[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11332_ _05377_ net590 _05607_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11263_ _05573_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13002_ clknet_leaf_81_clk _00460_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10214_ _04732_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__clkbuf_4
X_11194_ _05535_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__clkbuf_1
X_10145_ _04765_ rvsingle.dp.rf.rf\[28\]\[5\] _04930_ VGND VGND VPWR VPWR _04935_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10076_ _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__buf_2
XFILLER_0_89_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10978_ _05318_ rvsingle.dp.rf.rf\[31\]\[1\] _05419_ VGND VGND VPWR VPWR _05420_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12717_ clknet_leaf_45_clk _00175_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12648_ clknet_leaf_105_clk _00106_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12579_ clknet_leaf_121_clk _00037_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold306 rvsingle.dp.rf.rf\[28\]\[29\] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold317 rvsingle.dp.rf.rf\[23\]\[10\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 rvsingle.dp.rf.rf\[29\]\[29\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold339 rvsingle.dp.rf.rf\[2\]\[11\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _02473_ _02318_ _01580_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__o211a_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _04591_ _04600_ _04592_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__or3b_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _01137_ rvsingle.dp.rf.rf\[30\]\[15\] VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__nor2_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08672_ rvsingle.dp.rf.rf\[31\]\[14\] _01425_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07623_ _01828_ rvsingle.dp.rf.rf\[2\]\[4\] _01299_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_972 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07554_ _02469_ _02470_ _02472_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_75_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06505_ _01425_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07485_ rvsingle.dp.rf.rf\[9\]\[6\] _01561_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09224_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__buf_8
X_06436_ _01297_ rvsingle.dp.rf.rf\[31\]\[28\] _01303_ _01357_ VGND VGND VPWR VPWR
+ _01358_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06367_ _01085_ WriteData[29] _01180_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__a21o_1
X_09155_ _01210_ _04070_ _04074_ _01219_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08106_ rvsingle.dp.rf.rf\[19\]\[1\] _01124_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__or2b_1
X_09086_ rvsingle.dp.rf.rf\[25\]\[26\] _01943_ _01717_ _04005_ VGND VGND VPWR VPWR
+ _04006_ sky130_fd_sc_hd__o211a_1
X_06298_ _01215_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__buf_8
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08037_ rvsingle.dp.rf.rf\[7\]\[0\] _02929_ _02957_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09988_ _04801_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__clkbuf_4
X_08939_ rvsingle.dp.rf.rf\[1\]\[25\] _03778_ _01856_ VGND VGND VPWR VPWR _03860_
+ sky130_fd_sc_hd__o21ai_1
X_11950_ _05941_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10901_ _05374_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__clkbuf_1
X_11881_ _05728_ rvsingle.dp.rf.rf\[6\]\[2\] _05902_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__mux2_1
X_10832_ _05330_ net704 _05320_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10763_ _05288_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12502_ clknet_leaf_34_clk _00986_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10694_ _05250_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12433_ clknet_leaf_48_clk _00917_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12364_ clknet_leaf_52_clk _00848_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11315_ _05600_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12295_ _04718_ _06096_ _06097_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11246_ _05562_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11177_ _05523_ _05487_ _05524_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__o21ai_1
X_10128_ _04916_ _04918_ _04920_ _04922_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__and4_2
XFILLER_0_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10059_ _04861_ _04641_ _04743_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__mux2_2
XFILLER_0_54_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07270_ _02093_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06221_ Instr[24] VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__buf_8
XFILLER_0_72_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06152_ Instr[4] Instr[5] VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold103 rvsingle.dp.rf.rf\[3\]\[17\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold114 rvsingle.dp.rf.rf\[9\]\[13\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold125 rvsingle.dp.rf.rf\[11\]\[5\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
Xhold136 rvsingle.dp.rf.rf\[12\]\[0\] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold147 rvsingle.dp.rf.rf\[0\]\[0\] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 rvsingle.dp.rf.rf\[17\]\[14\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ Instr[7] VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__clkbuf_4
Xhold169 rvsingle.dp.rf.rf\[1\]\[19\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09842_ _04671_ _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__nand2_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _04606_ _04609_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__xnor2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _01900_ _01902_ _01721_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _02473_ _02318_ _01961_ _03644_ _01580_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _01425_ rvsingle.dp.rf.rf\[14\]\[14\] VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _01115_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__buf_6
XFILLER_0_139_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _03505_ _01335_ _01727_ _03506_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07537_ _01725_ rvsingle.dp.rf.rf\[22\]\[6\] _01198_ VGND VGND VPWR VPWR _02458_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_165_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07468_ _02383_ _01505_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__nand3_1
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09207_ _02907_ _02963_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__nor2_1
X_06419_ rvsingle.dp.rf.rf\[21\]\[29\] _01297_ _01310_ _01340_ VGND VGND VPWR VPWR
+ _01341_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_107_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07399_ _01551_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__clkbuf_8
X_09138_ _03983_ _04053_ _04056_ _04057_ _03982_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09069_ rvsingle.dp.rf.rf\[4\]\[26\] rvsingle.dp.rf.rf\[5\]\[26\] _01337_ VGND VGND
+ VPWR VPWR _03989_ sky130_fd_sc_hd__mux2_1
X_11100_ _05482_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__clkbuf_1
X_12080_ _05721_ _06007_ _06008_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__a21oi_1
Xhold670 rvsingle.dp.rf.rf\[21\]\[22\] VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 rvsingle.dp.rf.rf\[12\]\[1\] VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 rvsingle.dp.rf.rf\[17\]\[13\] VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _05448_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__clkbuf_1
X_12982_ clknet_leaf_31_clk _00440_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11933_ _05713_ net240 _05924_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _05716_ net661 _05885_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__mux2_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _05318_ net280 _05320_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__mux2_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11795_ _05856_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10746_ _05279_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10677_ _05241_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12416_ clknet_leaf_117_clk _00900_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13396_ clknet_leaf_21_clk _00824_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12347_ _06125_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12278_ _06088_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__clkbuf_1
X_11229_ _05300_ rvsingle.dp.rf.rf\[29\]\[22\] _05552_ VGND VGND VPWR VPWR _05554_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06770_ _01690_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__buf_8
XFILLER_0_78_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08440_ _01268_ rvsingle.dp.rf.rf\[22\]\[9\] _02059_ _03360_ VGND VGND VPWR VPWR
+ _03361_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_59_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08371_ rvsingle.dp.rf.rf\[9\]\[8\] _01424_ _01716_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07322_ _01269_ rvsingle.dp.rf.rf\[0\]\[16\] _02242_ _01497_ VGND VGND VPWR VPWR
+ _02243_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_105_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07253_ _01703_ _02173_ _01478_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06204_ _01127_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__buf_6
XFILLER_0_121_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07184_ rvsingle.dp.rf.rf\[25\]\[17\] _01847_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06135_ Instr[13] Instr[14] VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09825_ PC[19] PC[20] PC[21] _04657_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__and4_1
X_09756_ PC[20] _04582_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__xor2_1
X_06968_ _01885_ _01886_ _01888_ _01565_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__o211ai_1
X_08707_ _01618_ rvsingle.dp.rf.rf\[14\]\[14\] _01530_ VGND VGND VPWR VPWR _03628_
+ sky130_fd_sc_hd__o21a_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _04511_ _04518_ _04504_ _04528_ _04530_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__o311a_1
X_06899_ _01812_ _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__nand2_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _03553_ _03558_ _02527_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__nand3_2
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ rvsingle.dp.rf.rf\[12\]\[12\] rvsingle.dp.rf.rf\[13\]\[12\] rvsingle.dp.rf.rf\[14\]\[12\]
+ rvsingle.dp.rf.rf\[15\]\[12\] _02176_ _01696_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__mux4_2
XFILLER_0_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10600_ _05198_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11580_ _05750_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10531_ _04770_ net768 _05152_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13250_ clknet_leaf_121_clk _00708_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10462_ _04790_ rvsingle.dp.rf.rf\[24\]\[11\] _05110_ VGND VGND VPWR VPWR _05118_
+ sky130_fd_sc_hd__mux2_1
X_12201_ _05769_ _05770_ _06045_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13181_ clknet_leaf_139_clk _00639_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10393_ _05078_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12132_ _06036_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12063_ _05999_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__clkbuf_1
X_11014_ _04827_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__buf_2
XFILLER_0_95_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ clknet_leaf_108_clk _00423_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11916_ _04833_ net520 _05913_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__mux2_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ clknet_leaf_114_clk _00354_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11847_ _05862_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__buf_8
XFILLER_0_129_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _05398_ net547 _05845_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10729_ net58 VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13379_ clknet_leaf_124_clk _00807_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07940_ _02858_ _02859_ _02803_ _02860_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07871_ _01567_ rvsingle.dp.rf.rf\[20\]\[2\] _02791_ _02395_ VGND VGND VPWR VPWR
+ _02792_ sky130_fd_sc_hd__o211ai_1
X_09610_ _04438_ _04447_ _04448_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__and3_1
X_06822_ _01124_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__clkbuf_8
X_09541_ _04366_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__clkbuf_4
X_06753_ _01614_ rvsingle.dp.rf.rf\[18\]\[20\] VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__nor2_1
X_09472_ _04376_ VGND VGND VPWR VPWR MemWrite sky130_fd_sc_hd__buf_6
X_06684_ _01604_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__buf_8
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08423_ rvsingle.dp.rf.rf\[29\]\[9\] _01618_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__or2b_1
XFILLER_0_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08354_ rvsingle.dp.rf.rf\[21\]\[8\] _03258_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07305_ rvsingle.dp.rf.rf\[25\]\[16\] _02030_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08285_ _01567_ rvsingle.dp.rf.rf\[24\]\[10\] _01604_ VGND VGND VPWR VPWR _03206_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07236_ _01691_ rvsingle.dp.rf.rf\[6\]\[17\] VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07167_ _01915_ _02082_ _02087_ _01218_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_70_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07098_ _01595_ rvsingle.dp.rf.rf\[26\]\[18\] _01490_ VGND VGND VPWR VPWR _02019_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09808_ _04638_ _04452_ _04642_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[24\] sky130_fd_sc_hd__o21ai_1
X_09739_ _04573_ _04569_ _04571_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__o21ai_1
X_12750_ clknet_leaf_71_clk _00208_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _05391_ rvsingle.dp.rf.rf\[10\]\[14\] _05806_ VGND VGND VPWR VPWR _05810_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ clknet_leaf_95_clk _00139_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ net72 _05778_ _05739_ _05501_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11563_ _05741_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13302_ clknet_leaf_62_clk _00760_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10514_ Instr[11] _04724_ Instr[10] VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__or3b_1
XFILLER_0_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11494_ _05391_ net368 _05695_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13233_ clknet_leaf_27_clk _00691_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10445_ _05107_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13164_ clknet_leaf_84_clk _00622_ _00001_ VGND VGND VPWR VPWR PC[1] sky130_fd_sc_hd__dfrtp_4
X_10376_ _05070_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__clkbuf_1
X_12115_ _06027_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__clkbuf_1
X_13095_ clknet_leaf_101_clk _00553_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_12046_ _05344_ net537 _05983_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ clknet_leaf_22_clk _00406_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_170 _01707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ clknet_leaf_41_clk _00337_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_192 _02176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08070_ rvsingle.dp.rf.rf\[31\]\[1\] _01440_ _02162_ VGND VGND VPWR VPWR _02991_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07021_ _01222_ _01933_ _01935_ _01450_ _01941_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08972_ _01223_ _03883_ _03887_ _01189_ _03891_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__o311ai_4
X_07923_ _01335_ rvsingle.dp.rf.rf\[30\]\[2\] _01727_ _02843_ VGND VGND VPWR VPWR
+ _02844_ sky130_fd_sc_hd__o211ai_1
Xhold18 rvsingle.dp.rf.rf\[19\]\[10\] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 rvsingle.dp.rf.rf\[4\]\[31\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07854_ _01499_ rvsingle.dp.rf.rf\[30\]\[2\] VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__nor2_1
X_06805_ _01725_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__buf_8
X_07785_ _01607_ rvsingle.dp.rf.rf\[12\]\[3\] VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__nor2_1
X_09524_ _04301_ _04302_ VGND VGND VPWR VPWR DataAdr[11] sky130_fd_sc_hd__nand2_8
X_06736_ _01656_ rvsingle.dp.rf.rf\[24\]\[20\] VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09455_ _04274_ _04289_ _04361_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__nor3_1
X_06667_ _01587_ _01578_ _01486_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__a21o_1
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08406_ _01268_ rvsingle.dp.rf.rf\[14\]\[9\] _02059_ _03326_ VGND VGND VPWR VPWR
+ _03327_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09386_ _04294_ _04298_ _04136_ _04300_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__o211ai_4
X_06598_ _01103_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08337_ _01135_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08268_ rvsingle.dp.rf.rf\[5\]\[10\] _02005_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07219_ _01753_ rvsingle.dp.rf.rf\[4\]\[17\] VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08199_ _01828_ rvsingle.dp.rf.rf\[8\]\[11\] VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10230_ net30 _04978_ _04987_ _04985_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10161_ _04943_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__clkbuf_1
X_10092_ _04365_ _04889_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12802_ clknet_leaf_140_clk _00260_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10994_ _04781_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ clknet_leaf_143_clk _00191_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ clknet_leaf_33_clk _00122_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11615_ _05769_ _05770_ _05722_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12595_ clknet_leaf_35_clk _00053_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11546_ _05730_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11477_ _05496_ net627 _05684_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13216_ clknet_leaf_132_clk _00674_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10428_ _04909_ _04913_ _05059_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ clknet_leaf_142_clk _00605_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10359_ _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__clkbuf_4
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ clknet_leaf_24_clk _00536_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12029_ _05975_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__buf_8
XFILLER_0_79_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07570_ _01115_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__clkbuf_8
X_06521_ _01420_ rvsingle.dp.rf.rf\[22\]\[21\] VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09240_ _04153_ _04156_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_146_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06452_ _01219_ _01367_ _01373_ _01189_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09171_ rvsingle.dp.rf.rf\[29\]\[31\] _01090_ _01094_ _04090_ VGND VGND VPWR VPWR
+ _04091_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06383_ rvsingle.dp.rf.rf\[3\]\[29\] _01298_ _01304_ VGND VGND VPWR VPWR _01305_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08122_ _03019_ _01082_ _01152_ _03042_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__nand4_4
XFILLER_0_160_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08053_ _02969_ _02972_ _01207_ _02973_ _02438_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_24_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07004_ _01317_ _01914_ _01924_ _01247_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08955_ _03872_ _03873_ _03782_ _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__o211ai_1
X_07906_ _01420_ rvsingle.dp.rf.rf\[22\]\[2\] VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__nor2_1
X_08886_ _01451_ _03806_ _01445_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__a21oi_1
X_07837_ _01508_ rvsingle.dp.rf.rf\[13\]\[2\] _02757_ VGND VGND VPWR VPWR _02758_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07768_ rvsingle.dp.rf.rf\[24\]\[3\] rvsingle.dp.rf.rf\[25\]\[3\] rvsingle.dp.rf.rf\[26\]\[3\]
+ rvsingle.dp.rf.rf\[27\]\[3\] _02450_ _01708_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__mux4_1
X_09507_ _04390_ VGND VGND VPWR VPWR WriteData[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06719_ _01628_ _01633_ _01634_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_67_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07699_ _02614_ _02491_ _02619_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__nand3_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ _02751_ _02857_ _02862_ _03053_ _02577_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__a221o_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09369_ _01185_ _01405_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11400_ _05648_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__clkbuf_1
X_12380_ clknet_leaf_147_clk _00864_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_70 ReadData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 ReadData[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11331_ _05610_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_92 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11262_ _05377_ rvsingle.dp.rf.rf\[15\]\[4\] _05569_ VGND VGND VPWR VPWR _05573_
+ sky130_fd_sc_hd__mux2_1
X_13001_ clknet_leaf_97_clk _00459_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10213_ Instr[7] Instr[8] VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__nand2_2
X_11193_ _05534_ net752 _05528_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10144_ _04934_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10075_ _04875_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10977_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__buf_6
XFILLER_0_85_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12716_ clknet_leaf_50_clk _00174_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12647_ clknet_leaf_104_clk _00105_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12578_ clknet_leaf_128_clk _00036_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11529_ _05639_ net263 _05706_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold307 rvsingle.dp.rf.rf\[3\]\[23\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold318 rvsingle.dp.rf.rf\[21\]\[7\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 rvsingle.dp.rf.rf\[6\]\[10\] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _01853_ _03655_ _03660_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__nand3_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08671_ rvsingle.dp.rf.rf\[28\]\[14\] rvsingle.dp.rf.rf\[29\]\[14\] _01191_ VGND
+ VGND VPWR VPWR _03592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07622_ _01206_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__buf_6
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07553_ _02473_ _02102_ _02471_ _02431_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06504_ Instr[15] VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__buf_6
X_07484_ _01847_ rvsingle.dp.rf.rf\[8\]\[6\] _01551_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09223_ _04140_ _04141_ Instr[13] Instr[14] _02259_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__o2111a_4
X_06435_ _01337_ rvsingle.dp.rf.rf\[30\]\[28\] VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09154_ _01226_ _04071_ _04073_ _01232_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06366_ _01085_ WriteData[29] _01180_ _01184_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__a211o_2
XFILLER_0_115_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08105_ rvsingle.dp.rf.rf\[17\]\[1\] _01381_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09085_ _01432_ rvsingle.dp.rf.rf\[24\]\[26\] VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__or2_1
X_06297_ _01211_ _01214_ _01219_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08036_ _01240_ rvsingle.dp.rf.rf\[6\]\[0\] _01454_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09987_ _04800_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__clkbuf_4
X_08938_ _01127_ rvsingle.dp.rf.rf\[0\]\[25\] VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__nor2_1
X_08869_ _01117_ _03783_ _01682_ _03789_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_153_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10900_ _05318_ rvsingle.dp.rf.rf\[18\]\[1\] _05373_ VGND VGND VPWR VPWR _05374_
+ sky130_fd_sc_hd__mux2_1
X_11880_ _05903_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10831_ _04777_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10762_ _05209_ rvsingle.dp.rf.rf\[20\]\[13\] _05285_ VGND VGND VPWR VPWR _05288_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12501_ clknet_leaf_36_clk _00985_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10693_ _04808_ rvsingle.dp.rf.rf\[21\]\[14\] _05246_ VGND VGND VPWR VPWR _05250_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12432_ clknet_leaf_70_clk _00916_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12363_ clknet_leaf_88_clk _00847_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11314_ _05266_ net440 _05591_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12294_ _04728_ _04925_ net53 VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11245_ _05187_ net302 _05552_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11176_ _05364_ _05365_ _05487_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10127_ _04921_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__buf_2
X_10058_ DataAdr[24] ReadData[24] _04750_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06220_ _01119_ _01122_ _01143_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06151_ _01074_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold104 rvsingle.dp.rf.rf\[11\]\[15\] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 rvsingle.dp.rf.rf\[18\]\[0\] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 rvsingle.dp.rf.rf\[19\]\[14\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold137 rvsingle.dp.rf.rf\[17\]\[19\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold148 rvsingle.dp.rf.rf\[26\]\[0\] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09910_ _04735_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold159 rvsingle.dp.rf.rf\[17\]\[5\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09841_ _04617_ PC[28] VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__nand2_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _04607_ _04608_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__or2_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ rvsingle.dp.rf.rf\[17\]\[22\] _01424_ _01716_ _01904_ VGND VGND VPWR VPWR
+ _01905_ sky130_fd_sc_hd__o211ai_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _01962_ _01128_ _03620_ _03643_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08654_ rvsingle.dp.rf.rf\[12\]\[14\] rvsingle.dp.rf.rf\[13\]\[14\] _01828_ VGND
+ VGND VPWR VPWR _03575_ sky130_fd_sc_hd__mux2_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07605_ _01660_ _02522_ _02523_ _02351_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_77_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _01328_ rvsingle.dp.rf.rf\[20\]\[12\] VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07536_ rvsingle.dp.rf.rf\[21\]\[6\] _02271_ _02268_ VGND VGND VPWR VPWR _02457_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07467_ _01496_ _02384_ _02385_ _02323_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_146_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09206_ _01063_ _04122_ _04117_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06418_ _01337_ rvsingle.dp.rf.rf\[20\]\[29\] VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07398_ Instr[27] VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09137_ _03909_ _03827_ _03908_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__a21boi_1
X_06349_ _01113_ _01264_ _01266_ _01271_ _01118_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__o221a_1
XFILLER_0_161_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09068_ _03985_ _03986_ _03987_ _01310_ _01915_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08019_ _01725_ rvsingle.dp.rf.rf\[8\]\[0\] _01454_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__o21bai_1
Xhold660 rvsingle.dp.rf.rf\[7\]\[26\] VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold671 rvsingle.dp.rf.rf\[9\]\[4\] VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ _05304_ net637 _05443_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__mux2_1
Xhold682 rvsingle.dp.rf.rf\[12\]\[13\] VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 rvsingle.dp.rf.rf\[25\]\[27\] VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12981_ clknet_leaf_37_clk _00439_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11932_ _05930_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__clkbuf_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _05893_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__clkbuf_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__buf_8
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _05716_ net359 _05845_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10745_ _04765_ rvsingle.dp.rf.rf\[20\]\[5\] _05274_ VGND VGND VPWR VPWR _05279_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10676_ _04770_ rvsingle.dp.rf.rf\[21\]\[6\] _05235_ VGND VGND VPWR VPWR _05241_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12415_ clknet_leaf_2_clk _00899_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13395_ clknet_4_8_0_clk _00823_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12346_ _05132_ net401 _06121_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12277_ _05132_ net303 _06073_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11228_ _05553_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ _05515_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_807 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08370_ _01329_ rvsingle.dp.rf.rf\[8\]\[8\] VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07321_ rvsingle.dp.rf.rf\[1\]\[16\] _01595_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07252_ rvsingle.dp.rf.rf\[24\]\[17\] rvsingle.dp.rf.rf\[25\]\[17\] rvsingle.dp.rf.rf\[26\]\[17\]
+ rvsingle.dp.rf.rf\[27\]\[17\] _01469_ _01728_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06203_ _01126_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07183_ rvsingle.dp.rf.rf\[27\]\[17\] _01088_ _01626_ VGND VGND VPWR VPWR _02104_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06134_ PC[1] VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09824_ PC[16] PC[17] PC[18] _04656_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__and4_1
X_06967_ rvsingle.dp.rf.rf\[17\]\[22\] _01088_ _01092_ _01887_ VGND VGND VPWR VPWR
+ _01888_ sky130_fd_sc_hd__o211ai_1
X_09755_ _04589_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__xor2_1
X_08706_ _01677_ rvsingle.dp.rf.rf\[13\]\[14\] _03626_ VGND VGND VPWR VPWR _03627_
+ sky130_fd_sc_hd__o21ai_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09686_ _04527_ _04528_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__a21oi_1
X_06898_ _01703_ _01813_ _01818_ _01218_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__o211ai_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _03554_ _03555_ _02351_ _03557_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__o211ai_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _01207_ _03488_ _02447_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07519_ _01327_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__buf_6
X_08499_ _03418_ _03419_ _01564_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10530_ net88 _05155_ _05159_ _05157_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10461_ _05117_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12200_ net62 VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__inv_2
X_13180_ clknet_leaf_14_clk _00638_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10392_ _04802_ net818 _05071_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12131_ _05132_ net348 _06031_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12062_ _05132_ net409 _05994_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__mux2_1
Xhold490 rvsingle.dp.rf.rf\[30\]\[16\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11013_ _05438_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ clknet_leaf_110_clk _00422_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _05921_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__clkbuf_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ clknet_leaf_2_clk _00353_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _05884_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11777_ _05753_ _05847_ _05840_ net105 VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10728_ _05268_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10659_ _04909_ _04913_ _05191_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13378_ clknet_leaf_130_clk _00806_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12329_ _05344_ net490 _06110_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07870_ rvsingle.dp.rf.rf\[21\]\[2\] _01544_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__or2b_1
X_06821_ _01739_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__nand2_2
X_09540_ PC[2] VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__clkbuf_4
X_06752_ _01671_ _01672_ _01617_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__o21ai_1
X_09471_ _01067_ _02912_ _01071_ _01062_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__and4b_1
X_06683_ _01103_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_8
X_08422_ rvsingle.dp.rf.rf\[31\]\[9\] _01796_ _01660_ VGND VGND VPWR VPWR _03343_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08353_ _01763_ rvsingle.dp.rf.rf\[20\]\[8\] VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07304_ _02223_ _01257_ _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08284_ _01853_ _03199_ _03204_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__nand3_1
XFILLER_0_74_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07235_ rvsingle.dp.rf.rf\[4\]\[17\] rvsingle.dp.rf.rf\[5\]\[17\] _01417_ VGND VGND
+ VPWR VPWR _02156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07166_ _02083_ _02084_ _01703_ _02086_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_132_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07097_ rvsingle.dp.rf.rf\[25\]\[18\] _01861_ _01759_ VGND VGND VPWR VPWR _02018_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09807_ _04422_ _04423_ _04641_ _04427_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__o211ai_1
X_07999_ _01307_ _02916_ _02917_ _02919_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__o31ai_1
X_09738_ PC[19] _04577_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__xnor2_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09669_ Instr[13] _02912_ _04506_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _05809_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
X_12680_ clknet_leaf_105_clk _00138_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ net63 _05778_ _05738_ _05501_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__a22o_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11562_ _05740_ rvsingle.dp.rf.rf\[11\]\[8\] _05729_ VGND VGND VPWR VPWR _05741_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10513_ _04719_ _05143_ _05147_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__a21oi_1
X_13301_ clknet_leaf_29_clk _00759_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11493_ _05698_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13232_ clknet_leaf_53_clk _00690_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10444_ _04760_ net445 _05103_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13163_ clknet_leaf_74_clk _00621_ _00000_ VGND VGND VPWR VPWR PC[0] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10375_ _04760_ net586 _05065_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12114_ _05344_ net428 _06019_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__mux2_1
X_13094_ clknet_leaf_121_clk _00552_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_12045_ _05990_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12947_ clknet_leaf_34_clk _00405_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ clknet_leaf_52_clk _00336_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 _01707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_182 _01828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_193 _02288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11829_ _04795_ net696 _05874_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07020_ _01703_ _01936_ _01938_ _01940_ _01478_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_125_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08971_ _01209_ _03888_ _03890_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07922_ rvsingle.dp.rf.rf\[31\]\[2\] _01690_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__or2b_1
Xhold19 rvsingle.dp.rf.rf\[3\]\[7\] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _01377_ _02762_ _02773_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__nand3_4
X_06804_ _01190_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07784_ _01650_ rvsingle.dp.rf.rf\[14\]\[3\] _01647_ VGND VGND VPWR VPWR _02705_
+ sky130_fd_sc_hd__o21ai_1
X_06735_ _01561_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__buf_6
X_09523_ _04358_ VGND VGND VPWR VPWR DataAdr[6] sky130_fd_sc_hd__clkinv_8
XFILLER_0_78_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09454_ _04293_ _04307_ _04317_ _04360_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__nand4_2
X_06666_ _01580_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__buf_4
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08405_ rvsingle.dp.rf.rf\[15\]\[9\] _01492_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__or2b_1
X_09385_ _03227_ _04294_ _04299_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06597_ _01136_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__buf_8
XFILLER_0_164_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08336_ rvsingle.dp.rf.rf\[29\]\[8\] _01650_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__and2b_1
XFILLER_0_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08267_ _01780_ rvsingle.dp.rf.rf\[4\]\[10\] VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_140_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_140_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07218_ rvsingle.dp.rf.rf\[7\]\[17\] _01088_ _01626_ VGND VGND VPWR VPWR _02139_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08198_ rvsingle.dp.rf.rf\[11\]\[11\] _01295_ _01953_ VGND VGND VPWR VPWR _03119_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07149_ rvsingle.dp.rf.rf\[4\]\[18\] rvsingle.dp.rf.rf\[5\]\[18\] _01432_ VGND VGND
+ VPWR VPWR _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10160_ _04796_ net612 _04941_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__mux2_1
X_10091_ _04365_ _04679_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12801_ clknet_leaf_130_clk _00259_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10993_ _05427_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ clknet_leaf_147_clk _00190_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ clknet_leaf_7_clk _00121_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11614_ _04912_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12594_ clknet_leaf_39_clk _00052_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11545_ _05728_ rvsingle.dp.rf.rf\[11\]\[2\] _05729_ VGND VGND VPWR VPWR _05730_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_131_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_131_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11476_ _05689_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13215_ clknet_leaf_148_clk _00673_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10427_ net67 VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13146_ clknet_leaf_1_clk _00604_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10358_ _04919_ Instr[7] VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__nor2b_2
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ clknet_leaf_65_clk _00535_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10289_ net148 _05019_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12028_ _05982_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06520_ _01440_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06451_ _01232_ _01368_ _01370_ _01372_ _01224_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09170_ _01100_ rvsingle.dp.rf.rf\[28\]\[31\] VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06382_ _01195_ rvsingle.dp.rf.rf\[2\]\[29\] _01303_ VGND VGND VPWR VPWR _01304_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08121_ _03030_ _01145_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__nand3_4
XFILLER_0_161_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_122_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_122_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08052_ rvsingle.dp.rf.rf\[12\]\[1\] rvsingle.dp.rf.rf\[13\]\[1\] rvsingle.dp.rf.rf\[14\]\[1\]
+ rvsingle.dp.rf.rf\[15\]\[1\] _01903_ _01470_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07003_ _01316_ _01919_ _01923_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08954_ rvsingle.dp.rf.rf\[15\]\[25\] _03778_ _03874_ VGND VGND VPWR VPWR _03875_
+ sky130_fd_sc_hd__o21ai_1
X_07905_ _01315_ _02814_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__nand3_1
X_08885_ rvsingle.dp.rf.rf\[18\]\[24\] rvsingle.dp.rf.rf\[19\]\[24\] _01192_ VGND
+ VGND VPWR VPWR _03806_ sky130_fd_sc_hd__mux2_1
X_07836_ _01594_ rvsingle.dp.rf.rf\[12\]\[2\] _01258_ VGND VGND VPWR VPWR _02757_
+ sky130_fd_sc_hd__o21ba_1
X_07767_ _02302_ _02687_ _02447_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__o21ai_2
X_09506_ _04377_ _02346_ _02371_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__and3_1
X_06718_ _01612_ _01635_ _01636_ _01600_ _01638_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_149_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07698_ _01542_ _02615_ _02616_ _01502_ _02618_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__o311ai_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06649_ _01491_ _01560_ _01563_ _01565_ _01569_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__o311ai_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ _04340_ _04344_ net825 _01067_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__nand4_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09368_ _04278_ _04137_ _04281_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_164_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08319_ _01499_ rvsingle.dp.rf.rf\[10\]\[8\] VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_113_clk sky130_fd_sc_hd__clkbuf_16
X_09299_ _04213_ _04214_ _03765_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__or3_1
XANTENNA_60 ReadData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_71 ReadData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ _05531_ rvsingle.dp.rf.rf\[14\]\[3\] _05607_ VGND VGND VPWR VPWR _05610_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_82 ReadData[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_93 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11261_ _05572_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13000_ clknet_leaf_105_clk _00458_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10212_ _04719_ _04969_ _04974_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11192_ _04764_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__buf_2
X_10143_ _04760_ net774 _04930_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10074_ _04364_ _04873_ _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10976_ _04927_ _04928_ _05417_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__or3_2
X_12715_ clknet_leaf_86_clk _00173_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12646_ clknet_leaf_113_clk _00104_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_104_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_104_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12577_ clknet_leaf_130_clk _00035_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11528_ _05717_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold308 rvsingle.dp.rf.rf\[25\]\[24\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold319 rvsingle.dp.rf.rf\[1\]\[25\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11459_ net59 VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13129_ clknet_leaf_92_clk _00587_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08670_ rvsingle.dp.rf.rf\[24\]\[14\] rvsingle.dp.rf.rf\[25\]\[14\] rvsingle.dp.rf.rf\[26\]\[14\]
+ rvsingle.dp.rf.rf\[27\]\[14\] _01426_ _01433_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__mux4_1
X_07621_ rvsingle.dp.rf.rf\[4\]\[4\] rvsingle.dp.rf.rf\[5\]\[4\] rvsingle.dp.rf.rf\[6\]\[4\]
+ rvsingle.dp.rf.rf\[7\]\[4\] _01416_ _01300_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__mux4_1
X_07552_ _01064_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_996 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06503_ _01423_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__clkbuf_8
X_07483_ _01763_ rvsingle.dp.rf.rf\[10\]\[6\] _02031_ _02403_ VGND VGND VPWR VPWR
+ _02404_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06434_ rvsingle.dp.rf.rf\[28\]\[28\] rvsingle.dp.rf.rf\[29\]\[28\] _01194_ VGND
+ VGND VPWR VPWR _01356_ sky130_fd_sc_hd__mux2_1
X_09222_ _01072_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09153_ rvsingle.dp.rf.rf\[1\]\[31\] _01298_ _01311_ _04072_ VGND VGND VPWR VPWR
+ _04073_ sky130_fd_sc_hd__o211a_1
X_06365_ _01147_ _01273_ _01287_ _01154_ VGND VGND VPWR VPWR WriteData[29] sky130_fd_sc_hd__o211a_4
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08104_ _01602_ rvsingle.dp.rf.rf\[16\]\[1\] VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09084_ rvsingle.dp.rf.rf\[26\]\[26\] rvsingle.dp.rf.rf\[27\]\[26\] _01193_ VGND
+ VGND VPWR VPWR _04004_ sky130_fd_sc_hd__mux2_1
X_06296_ _01218_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08035_ rvsingle.dp.rf.rf\[5\]\[0\] _01423_ _01307_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09986_ _04799_ _04524_ _04364_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__mux2_4
XFILLER_0_110_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08937_ rvsingle.dp.rf.rf\[3\]\[25\] _03857_ _03840_ VGND VGND VPWR VPWR _03858_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08868_ _01512_ _03784_ _03786_ _03788_ _01506_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07819_ rvsingle.dp.rf.rf\[17\]\[3\] _01544_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__and2b_1
X_08799_ rvsingle.dp.rf.rf\[4\]\[15\] rvsingle.dp.rf.rf\[5\]\[15\] rvsingle.dp.rf.rf\[6\]\[15\]
+ rvsingle.dp.rf.rf\[7\]\[15\] _01335_ _01244_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__mux4_1
X_10830_ _05329_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10761_ _05287_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12500_ clknet_leaf_21_clk _00984_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10692_ _05249_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12431_ clknet_leaf_39_clk _00915_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12362_ _06132_ _06096_ _06133_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11313_ _05599_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__clkbuf_1
X_12293_ _04916_ _04918_ _04728_ _04922_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__and4_2
XFILLER_0_132_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11244_ _05561_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11175_ net46 VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__inv_2
X_10126_ _02909_ _02910_ _02799_ _04724_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__o31a_2
XFILLER_0_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10057_ _04860_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10959_ _05407_ net746 _05401_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12629_ clknet_leaf_36_clk _00087_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06150_ _01073_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__buf_4
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold105 rvsingle.dp.rf.rf\[7\]\[19\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold116 rvsingle.dp.rf.rf\[4\]\[0\] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 rvsingle.dp.rf.rf\[21\]\[0\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold138 rvsingle.dp.rf.rf\[3\]\[3\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 rvsingle.dp.rf.rf\[8\]\[0\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _04617_ PC[28] VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__or2_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _04590_ PC[22] VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__nor2_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _01903_ rvsingle.dp.rf.rf\[16\]\[22\] VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__or2_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _01377_ _03631_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__nand3_4
X_08653_ rvsingle.dp.rf.rf\[8\]\[14\] rvsingle.dp.rf.rf\[9\]\[14\] rvsingle.dp.rf.rf\[10\]\[14\]
+ rvsingle.dp.rf.rf\[11\]\[14\] _01730_ _01953_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07604_ rvsingle.dp.rf.rf\[27\]\[4\] _01487_ _02524_ VGND VGND VPWR VPWR _02525_
+ sky130_fd_sc_hd__o21ai_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ rvsingle.dp.rf.rf\[21\]\[12\] VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07535_ _01420_ rvsingle.dp.rf.rf\[20\]\[6\] VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07466_ _02379_ rvsingle.dp.rf.rf\[29\]\[6\] _02386_ VGND VGND VPWR VPWR _02387_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06417_ rvsingle.dp.rf.rf\[16\]\[29\] rvsingle.dp.rf.rf\[17\]\[29\] rvsingle.dp.rf.rf\[18\]\[29\]
+ rvsingle.dp.rf.rf\[19\]\[29\] _01338_ _01303_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09205_ _02962_ _02964_ _02965_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__and3b_1
X_07397_ _01074_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__buf_8
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06348_ _01261_ _01270_ _01133_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__a21o_1
X_09136_ _03984_ _04055_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__nor2_2
XFILLER_0_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09067_ rvsingle.dp.rf.rf\[0\]\[26\] rvsingle.dp.rf.rf\[1\]\[26\] _01337_ VGND VGND
+ VPWR VPWR _03987_ sky130_fd_sc_hd__mux2_1
X_06279_ _01201_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08018_ _02926_ _02938_ _01187_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__nand3_2
XFILLER_0_102_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold650 rvsingle.dp.rf.rf\[21\]\[5\] VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold661 rvsingle.dp.rf.rf\[23\]\[29\] VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 rvsingle.dp.rf.rf\[22\]\[4\] VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold683 rvsingle.dp.rf.rf\[21\]\[8\] VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold694 rvsingle.dp.rf.rf\[22\]\[10\] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09969_ _04785_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__clkbuf_4
X_12980_ clknet_leaf_22_clk _00438_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11931_ _04876_ net579 _05924_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11862_ _05763_ net235 _05885_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__mux2_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10813_ _04722_ _04723_ _04965_ _05063_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__or4_4
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _05855_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__clkbuf_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10744_ _05278_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10675_ _05240_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12414_ clknet_leaf_2_clk _00898_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13394_ clknet_leaf_40_clk _00822_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12345_ _06124_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12276_ _06087_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11227_ _05400_ rvsingle.dp.rf.rf\[29\]\[21\] _05552_ VGND VGND VPWR VPWR _05553_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11158_ _05300_ net220 _05511_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__mux2_1
X_10109_ _04905_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
X_11089_ _05177_ _05471_ _05463_ net208 VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_136_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07320_ _01488_ rvsingle.dp.rf.rf\[3\]\[16\] _01491_ _02240_ VGND VGND VPWR VPWR
+ _02241_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07251_ _02169_ _01717_ _01722_ _02171_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06202_ _01125_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__buf_6
XFILLER_0_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07182_ _01666_ rvsingle.dp.rf.rf\[26\]\[17\] VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09823_ PC[13] PC[14] PC[15] _04655_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__and4_1
X_09754_ _04591_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__or2b_1
X_06966_ _01642_ rvsingle.dp.rf.rf\[16\]\[22\] VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__or2_1
X_08705_ _01255_ rvsingle.dp.rf.rf\[12\]\[14\] _01551_ VGND VGND VPWR VPWR _03626_
+ sky130_fd_sc_hd__o21ba_1
X_09685_ PC[14] _04529_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__xnor2_1
X_06897_ _01814_ _01815_ _01816_ _01817_ _01445_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__o221ai_2
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ rvsingle.dp.rf.rf\[27\]\[12\] _01487_ _03556_ VGND VGND VPWR VPWR _03557_
+ sky130_fd_sc_hd__o21ai_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08567_ rvsingle.dp.rf.rf\[4\]\[12\] rvsingle.dp.rf.rf\[5\]\[12\] rvsingle.dp.rf.rf\[6\]\[12\]
+ rvsingle.dp.rf.rf\[7\]\[12\] _02450_ _01708_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07518_ _01207_ _02437_ _02438_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_147_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08498_ rvsingle.dp.rf.rf\[17\]\[13\] _01498_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07449_ _02360_ _02363_ _02364_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10460_ _04786_ rvsingle.dp.rf.rf\[24\]\[10\] _05110_ VGND VGND VPWR VPWR _05117_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09119_ _01666_ rvsingle.dp.rf.rf\[18\]\[26\] _01626_ VGND VGND VPWR VPWR _04039_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10391_ _05077_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12130_ _06035_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12061_ _05998_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold480 rvsingle.dp.rf.rf\[25\]\[15\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 rvsingle.dp.rf.rf\[18\]\[7\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ _04824_ rvsingle.dp.rf.rf\[31\]\[17\] _05431_ VGND VGND VPWR VPWR _05438_
+ sky130_fd_sc_hd__mux2_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12963_ clknet_leaf_116_clk _00421_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_84_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _05173_ net414 _05913_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ clknet_leaf_150_clk _00352_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11845_ _04839_ net505 _05874_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__mux2_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _05848_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__clkbuf_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10727_ _05187_ net326 _05257_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10658_ net40 VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13377_ clknet_leaf_125_clk _00805_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10589_ net34 _05191_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12328_ _06115_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12259_ _05472_ _05847_ _06077_ net170 VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06820_ _01740_ _01685_ _01737_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__o21bai_1
X_06751_ rvsingle.dp.rf.rf\[21\]\[20\] _01558_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_75_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
X_06682_ _01602_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__buf_8
X_09470_ _04375_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08421_ _01603_ rvsingle.dp.rf.rf\[30\]\[9\] VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08352_ _01531_ _03269_ _03270_ _01131_ _03272_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_47_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07303_ _01098_ rvsingle.dp.rf.rf\[26\]\[16\] _01260_ VGND VGND VPWR VPWR _02224_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08283_ _01092_ _03200_ _03201_ _01511_ _03203_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07234_ _01703_ _02154_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07165_ rvsingle.dp.rf.rf\[23\]\[18\] _01943_ _02085_ VGND VGND VPWR VPWR _02086_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07096_ _01383_ rvsingle.dp.rf.rf\[24\]\[18\] VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09806_ _04639_ _04640_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__nor2_2
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07998_ _01423_ rvsingle.dp.rf.rf\[25\]\[0\] _02918_ VGND VGND VPWR VPWR _02919_
+ sky130_fd_sc_hd__o21ai_1
X_09737_ _01189_ _02912_ _01175_ _04507_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06949_ _01082_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_66_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
X_09668_ _04512_ _04453_ _04514_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[12\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _01382_ rvsingle.dp.rf.rf\[22\]\[12\] _02337_ VGND VGND VPWR VPWR _03540_
+ sky130_fd_sc_hd__o21ai_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _04449_ _04450_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__xnor2_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ net196 _05779_ _05736_ _05501_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11561_ _04777_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__buf_2
XFILLER_0_108_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13300_ clknet_leaf_58_clk _00758_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10512_ _05145_ _05146_ net1 VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__a21oi_1
X_11492_ _04801_ net682 _05695_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13231_ clknet_leaf_45_clk _00689_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10443_ _05106_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13162_ clknet_leaf_82_clk _00620_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10374_ _04984_ _05068_ _05069_ _05065_ net5 VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12113_ _06026_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13093_ clknet_leaf_110_clk _00551_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12044_ _04813_ net381 _05983_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_57_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ clknet_leaf_41_clk _00404_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ clknet_leaf_43_clk _00335_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_150 _01611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _01711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11828_ _05875_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_183 _01877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 _03139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11759_ _05840_ net92 _05739_ _05841_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08970_ _01231_ _03889_ _01223_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__o21a_1
X_07921_ rvsingle.dp.rf.rf\[29\]\[2\] _01687_ _02268_ _02841_ VGND VGND VPWR VPWR
+ _02842_ sky130_fd_sc_hd__o211ai_1
X_07852_ _02765_ _02767_ _02364_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__o211ai_2
X_06803_ _01722_ _01723_ _01218_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__o21ai_1
X_07783_ rvsingle.dp.rf.rf\[15\]\[3\] _01566_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_48_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09522_ _04354_ VGND VGND VPWR VPWR DataAdr[5] sky130_fd_sc_hd__inv_6
X_06734_ _01654_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__clkbuf_8
X_09453_ DataAdr[12] net819 DataAdr[9] _04359_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__nor4_1
X_06665_ _01480_ _01453_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08404_ rvsingle.dp.rf.rf\[13\]\[9\] _01743_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09384_ _04296_ _04297_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__nand2_1
X_06596_ _01495_ _01504_ _01506_ _01516_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_93_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08335_ _01878_ rvsingle.dp.rf.rf\[28\]\[8\] VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08266_ _01518_ rvsingle.dp.rf.rf\[2\]\[10\] _02320_ _03186_ VGND VGND VPWR VPWR
+ _03187_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07217_ _01666_ rvsingle.dp.rf.rf\[6\]\[17\] VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08197_ _01726_ rvsingle.dp.rf.rf\[10\]\[11\] VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07148_ rvsingle.dp.rf.rf\[0\]\[18\] rvsingle.dp.rf.rf\[1\]\[18\] rvsingle.dp.rf.rf\[2\]\[18\]
+ rvsingle.dp.rf.rf\[3\]\[18\] _01193_ _01451_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__mux4_2
XFILLER_0_113_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07079_ rvsingle.dp.rf.rf\[3\]\[19\] _01255_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10090_ _02908_ DataAdr[28] _04888_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
X_12800_ clknet_leaf_120_clk _00258_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10992_ _05330_ net737 _05419_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__mux2_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ clknet_leaf_141_clk _00189_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ clknet_leaf_33_clk _00120_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _04908_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__buf_2
XFILLER_0_108_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12593_ clknet_leaf_49_clk _00051_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11544_ _05725_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__buf_8
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11475_ _05534_ rvsingle.dp.rf.rf\[12\]\[5\] _05684_ VGND VGND VPWR VPWR _05689_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13214_ clknet_leaf_148_clk _00672_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10426_ _05094_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13145_ clknet_leaf_9_clk _00603_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10357_ _05055_ _05019_ _05056_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__o21ai_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ clknet_leaf_21_clk _00534_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10288_ _04721_ _04728_ _04966_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__and3_2
X_12027_ _04769_ net390 _05976_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12929_ clknet_leaf_117_clk _00387_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_06450_ _01202_ _01371_ _01209_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06381_ _01302_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08120_ _03035_ _01115_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__nand3_1
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08051_ _01460_ _02971_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07002_ _01915_ _01920_ _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08953_ _01666_ rvsingle.dp.rf.rf\[14\]\[25\] _01612_ VGND VGND VPWR VPWR _03874_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07904_ _01229_ _02819_ _02824_ _01217_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_138_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08884_ rvsingle.dp.rf.rf\[17\]\[24\] _01296_ _01717_ _03804_ VGND VGND VPWR VPWR
+ _03805_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_99_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07835_ _02752_ _02753_ _01131_ _02755_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07766_ rvsingle.dp.rf.rf\[16\]\[3\] rvsingle.dp.rf.rf\[17\]\[3\] rvsingle.dp.rf.rf\[18\]\[3\]
+ rvsingle.dp.rf.rf\[19\]\[3\] _01328_ _01455_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09505_ _04389_ VGND VGND VPWR VPWR WriteData[8] sky130_fd_sc_hd__inv_2
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06717_ _01619_ rvsingle.dp.rf.rf\[2\]\[20\] _01620_ _01637_ VGND VGND VPWR VPWR
+ _01638_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_52_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07697_ _01645_ rvsingle.dp.rf.rf\[13\]\[5\] _02617_ VGND VGND VPWR VPWR _02618_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _04341_ _04342_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__a21oi_4
X_06648_ _01559_ rvsingle.dp.rf.rf\[2\]\[21\] _01260_ _01568_ VGND VGND VPWR VPWR
+ _01569_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_149_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09367_ _04282_ _04122_ _04141_ _02012_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__and4bb_1
X_06579_ _01499_ rvsingle.dp.rf.rf\[24\]\[21\] VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08318_ rvsingle.dp.rf.rf\[9\]\[8\] _01539_ _01542_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__o21ai_1
X_09298_ _02098_ _02100_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__nand2_2
XANTENNA_50 ReadData[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_61 ReadData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 ReadData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_83 ReadData[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08249_ _03154_ _03169_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_94 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11260_ _05531_ rvsingle.dp.rf.rf\[15\]\[3\] _05569_ VGND VGND VPWR VPWR _05572_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10211_ _04970_ _04973_ net7 VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11191_ _05533_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__clkbuf_1
X_10142_ _04933_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__clkbuf_1
X_10073_ _04660_ _01080_ _04661_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__or3b_2
XFILLER_0_98_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10975_ _04975_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__buf_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ clknet_leaf_95_clk _00172_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12645_ clknet_leaf_115_clk _00103_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12576_ clknet_leaf_120_clk _00034_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11527_ _05716_ net222 _05706_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold309 rvsingle.dp.rf.rf\[12\]\[28\] VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11458_ _05678_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10409_ _04853_ net234 _05082_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__mux2_1
X_11389_ net71 VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__inv_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ clknet_leaf_101_clk _00586_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ clknet_leaf_125_clk _00517_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07620_ _01711_ _02535_ _02540_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07551_ _02471_ _02431_ _01591_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_159_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06502_ _01293_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_8
X_07482_ rvsingle.dp.rf.rf\[11\]\[6\] _01877_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09221_ _02260_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__clkbuf_4
X_06433_ rvsingle.dp.rf.rf\[24\]\[28\] rvsingle.dp.rf.rf\[25\]\[28\] rvsingle.dp.rf.rf\[26\]\[28\]
+ rvsingle.dp.rf.rf\[27\]\[28\] _01338_ _01202_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09152_ _01195_ rvsingle.dp.rf.rf\[0\]\[31\] VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__or2_1
X_06364_ _01118_ _01275_ _01279_ _01286_ _01147_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_17_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08103_ _01880_ _03020_ _03021_ _01110_ _03023_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_127_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09083_ rvsingle.dp.rf.rf\[28\]\[26\] rvsingle.dp.rf.rf\[29\]\[26\] rvsingle.dp.rf.rf\[30\]\[26\]
+ rvsingle.dp.rf.rf\[31\]\[26\] _01330_ _01302_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_886 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06295_ _01217_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__buf_6
X_08034_ _02176_ rvsingle.dp.rf.rf\[4\]\[0\] VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold810 rvsingle.dp.rf.rf\[14\]\[21\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09985_ ReadData[13] _04713_ _04245_ _04798_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08936_ _01646_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__clkbuf_4
X_08867_ _01491_ _03787_ _01768_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07818_ _01650_ rvsingle.dp.rf.rf\[16\]\[3\] VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__nor2_1
X_08798_ _01461_ _03714_ _03718_ _01447_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_98_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07749_ _01828_ rvsingle.dp.rf.rf\[2\]\[3\] VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10760_ _05207_ rvsingle.dp.rf.rf\[20\]\[12\] _05285_ VGND VGND VPWR VPWR _05287_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09419_ _04327_ _04328_ _04329_ VGND VGND VPWR VPWR DataAdr[9] sky130_fd_sc_hd__o21ai_4
XFILLER_0_66_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10691_ _05209_ rvsingle.dp.rf.rf\[21\]\[13\] _05246_ VGND VGND VPWR VPWR _05249_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12430_ clknet_leaf_67_clk _00914_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12361_ _04908_ _04912_ _06096_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11312_ _05359_ net449 _05591_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12292_ _06094_ _06070_ _06095_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11243_ _05266_ net328 _05552_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__mux2_1
X_11174_ _05522_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10125_ _04737_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__nor2_4
X_10056_ _04859_ net582 _04847_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10958_ _04875_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__buf_2
XFILLER_0_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10889_ _04912_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__buf_2
XFILLER_0_26_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12628_ clknet_leaf_59_clk _00086_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12559_ clknet_leaf_57_clk _01043_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold106 rvsingle.dp.rf.rf\[27\]\[6\] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 rvsingle.dp.rf.rf\[7\]\[6\] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold128 rvsingle.dp.rf.rf\[5\]\[13\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold139 rvsingle.dp.rf.rf\[9\]\[14\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _04590_ PC[22] VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__and2_1
X_06982_ _01327_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__buf_8
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _01853_ _03636_ _03641_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__nand3_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ net820 _03483_ _03565_ _03567_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__o2111ai_4
X_07603_ _01136_ rvsingle.dp.rf.rf\[26\]\[4\] _01551_ VGND VGND VPWR VPWR _02524_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08583_ rvsingle.dp.rf.rf\[16\]\[12\] rvsingle.dp.rf.rf\[17\]\[12\] rvsingle.dp.rf.rf\[18\]\[12\]
+ rvsingle.dp.rf.rf\[19\]\[12\] _01730_ _01808_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07534_ rvsingle.dp.rf.rf\[16\]\[6\] rvsingle.dp.rf.rf\[17\]\[6\] rvsingle.dp.rf.rf\[18\]\[6\]
+ rvsingle.dp.rf.rf\[19\]\[6\] _01462_ _01727_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07465_ _01779_ rvsingle.dp.rf.rf\[28\]\[6\] _01610_ VGND VGND VPWR VPWR _02386_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09204_ _04121_ _04122_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__or2_4
XFILLER_0_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06416_ _01337_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__buf_4
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07396_ _01188_ _02293_ _02316_ _01246_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09135_ _04053_ _04054_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__or2_2
XFILLER_0_162_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06347_ rvsingle.dp.rf.rf\[14\]\[29\] rvsingle.dp.rf.rf\[15\]\[29\] _01269_ VGND
+ VGND VPWR VPWR _01270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09066_ _01337_ rvsingle.dp.rf.rf\[2\]\[26\] VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06278_ _01200_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08017_ _01217_ _02932_ _02937_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 rvsingle.dp.rf.rf\[13\]\[11\] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold651 rvsingle.dp.rf.rf\[30\]\[19\] VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold662 rvsingle.dp.rf.rf\[22\]\[27\] VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold673 rvsingle.dp.rf.rf\[16\]\[19\] VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 rvsingle.dp.rf.rf\[3\]\[1\] VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 rvsingle.dp.rf.rf\[12\]\[19\] VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__dlygate4sd3_1
X_09968_ _04784_ _04479_ _04743_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__mux2_4
X_08919_ _01531_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__clkbuf_4
X_09899_ _04725_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__buf_4
X_11930_ _05929_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _05892_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__clkbuf_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _04735_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _05763_ net277 _05845_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10743_ _04760_ net807 _05274_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10674_ _04765_ net650 _05235_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12413_ clknet_leaf_143_clk _00897_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13393_ clknet_leaf_48_clk _00821_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12344_ _04858_ net226 _06121_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12275_ _04858_ net596 _06073_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11226_ _05527_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__buf_6
X_11157_ _05514_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10108_ _04904_ net233 _04847_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__mux2_1
X_11088_ _05478_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__clkbuf_1
X_10039_ _04365_ _04843_ _04844_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_59_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07250_ _01688_ rvsingle.dp.rf.rf\[31\]\[17\] _01301_ _02170_ VGND VGND VPWR VPWR
+ _02171_ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06201_ _01124_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_170_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07181_ _01074_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__buf_6
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09822_ PC[10] PC[11] PC[12] _04475_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09753_ Instr[31] PC[20] VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__or2_1
X_06965_ rvsingle.dp.rf.rf\[19\]\[22\] _01088_ _01626_ VGND VGND VPWR VPWR _01886_
+ sky130_fd_sc_hd__o21ai_1
X_08704_ _03621_ _03622_ _03624_ _02483_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__o211ai_1
X_09684_ Instr[14] _04505_ _04506_ _04507_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__a31o_1
X_06896_ rvsingle.dp.rf.rf\[7\]\[23\] _01688_ _01456_ VGND VGND VPWR VPWR _01817_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08635_ _01613_ rvsingle.dp.rf.rf\[26\]\[12\] _01551_ VGND VGND VPWR VPWR _03556_
+ sky130_fd_sc_hd__o21a_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _03484_ _01309_ _01229_ _03486_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_166_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07517_ _01215_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__clkbuf_8
X_08497_ _01769_ rvsingle.dp.rf.rf\[16\]\[13\] _01519_ VGND VGND VPWR VPWR _03418_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_147_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07448_ _01552_ _02365_ _02366_ _02329_ _02368_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_146_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07379_ _02295_ _02296_ _01721_ _02299_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_33_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09118_ rvsingle.dp.rf.rf\[17\]\[26\] _03839_ _01856_ VGND VGND VPWR VPWR _04038_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10390_ _04796_ net764 _05071_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09049_ _01138_ rvsingle.dp.rf.rf\[8\]\[27\] VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12060_ _05757_ net242 _05994_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold470 rvsingle.dp.rf.rf\[8\]\[19\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 rvsingle.dp.rf.rf\[30\]\[5\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ _05437_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__clkbuf_1
Xhold492 rvsingle.dp.rf.rf\[6\]\[14\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ clknet_leaf_141_clk _00420_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _05920_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__clkbuf_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ clknet_leaf_142_clk _00351_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _05883_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11775_ _05173_ net714 _05845_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _05267_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10657_ _05229_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13376_ clknet_leaf_120_clk _00804_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10588_ _04918_ _04728_ _04922_ _04916_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__and4b_2
XFILLER_0_106_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12327_ _04813_ net688 _06110_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12258_ _06081_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__clkbuf_1
X_11209_ _05543_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__clkbuf_1
X_12189_ _04982_ _04983_ _04981_ _05003_ net388 VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__o41a_1
XFILLER_0_76_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06750_ _01137_ rvsingle.dp.rf.rf\[20\]\[20\] _01611_ VGND VGND VPWR VPWR _01671_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_92_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06681_ _01135_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__buf_6
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08420_ _01593_ _03329_ _03340_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__nand3_2
XFILLER_0_86_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08351_ _01545_ rvsingle.dp.rf.rf\[18\]\[8\] _02031_ _03271_ VGND VGND VPWR VPWR
+ _03272_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_86_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07302_ rvsingle.dp.rf.rf\[27\]\[16\] VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08282_ _02481_ rvsingle.dp.rf.rf\[21\]\[10\] _03202_ VGND VGND VPWR VPWR _03203_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07233_ rvsingle.dp.rf.rf\[0\]\[17\] rvsingle.dp.rf.rf\[1\]\[17\] rvsingle.dp.rf.rf\[2\]\[17\]
+ rvsingle.dp.rf.rf\[3\]\[17\] _01726_ _01728_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07164_ _01432_ rvsingle.dp.rf.rf\[22\]\[18\] _01728_ VGND VGND VPWR VPWR _02085_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07095_ _01248_ _01942_ _01958_ _02012_ _02014_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__a32o_1
XFILLER_0_100_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09805_ PC[23] _04612_ PC[24] VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__a21oi_1
X_07997_ _01425_ rvsingle.dp.rf.rf\[24\]\[0\] _01197_ VGND VGND VPWR VPWR _02918_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06948_ _01846_ _01854_ _01859_ _01868_ _01378_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__o221ai_4
X_09736_ _04574_ _04453_ _04576_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[18\] sky130_fd_sc_hd__o21ai_1
X_09667_ _04454_ _04455_ _04513_ _04459_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__o211ai_1
X_06879_ _01668_ _01794_ _01795_ _01617_ _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_96_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _03505_ _01603_ _01660_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__a211oi_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ Instr[26] PC[6] _04442_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__a21oi_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _01240_ rvsingle.dp.rf.rf\[14\]\[13\] _01454_ VGND VGND VPWR VPWR _03470_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11560_ net11 _05726_ _05739_ _05737_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10511_ _05142_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11491_ _05697_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13230_ clknet_leaf_54_clk _00688_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10442_ _04755_ net731 _05103_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_973 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13161_ clknet_leaf_95_clk _00619_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10373_ _05060_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__buf_6
XFILLER_0_131_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12112_ _04813_ net532 _06019_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__mux2_1
X_13092_ clknet_leaf_101_clk _00550_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12043_ _05989_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ clknet_leaf_42_clk _00403_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ clknet_leaf_51_clk _00334_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_140 _01567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _01611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_162 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 _01726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 _01877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11827_ _05744_ net780 _05874_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__mux2_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _03139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _05840_ net117 _05738_ _05841_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10709_ _05258_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11689_ _05803_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13359_ clknet_leaf_66_clk _00787_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07920_ _01690_ rvsingle.dp.rf.rf\[28\]\[2\] VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__or2_1
X_07851_ _01490_ _02768_ _02769_ _01111_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__o311ai_2
X_06802_ rvsingle.dp.rf.rf\[20\]\[20\] rvsingle.dp.rf.rf\[21\]\[20\] rvsingle.dp.rf.rf\[22\]\[20\]
+ rvsingle.dp.rf.rf\[23\]\[20\] _01192_ _01244_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__mux4_1
X_07782_ _02699_ _02700_ _01564_ _02702_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__o211ai_1
X_09521_ _04344_ VGND VGND VPWR VPWR DataAdr[2] sky130_fd_sc_hd__inv_6
X_06733_ _01610_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ DataAdr[8] _04349_ _04354_ _04358_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_148_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06664_ _01153_ _01536_ _01577_ _01482_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__a41o_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08403_ _01268_ rvsingle.dp.rf.rf\[12\]\[9\] VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09383_ _04296_ _04297_ _03227_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__a21boi_2
X_06595_ _01507_ _01510_ _01512_ _01515_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08334_ _01593_ _03243_ _03254_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__nand3_4
XFILLER_0_129_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08265_ rvsingle.dp.rf.rf\[3\]\[10\] _01561_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07216_ _02128_ _02131_ _01526_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08196_ rvsingle.dp.rf.rf\[12\]\[11\] rvsingle.dp.rf.rf\[13\]\[11\] rvsingle.dp.rf.rf\[14\]\[11\]
+ rvsingle.dp.rf.rf\[15\]\[11\] _01416_ _01300_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__mux4_2
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07147_ _01587_ _02067_ _01486_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07078_ rvsingle.dp.rf.rf\[1\]\[19\] _01847_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_870 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09719_ _04547_ _04552_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__nor2_1
X_10991_ _05426_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__clkbuf_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ clknet_leaf_4_clk _00188_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ clknet_leaf_36_clk _00119_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11612_ net55 VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__inv_2
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ clknet_leaf_71_clk _00050_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11543_ _04746_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11474_ _05688_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13213_ clknet_leaf_139_clk _00671_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10425_ _04904_ net371 _05082_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13144_ clknet_leaf_28_clk _00602_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10356_ _04909_ _04913_ _05019_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ clknet_leaf_29_clk _00533_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10287_ _05017_ _04969_ _05018_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__o21ai_1
X_12026_ _05981_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12928_ clknet_leaf_116_clk _00386_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ clknet_leaf_142_clk _00317_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06380_ _01301_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__buf_4
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08050_ rvsingle.dp.rf.rf\[9\]\[1\] _02271_ _02268_ _02970_ VGND VGND VPWR VPWR _02971_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_109_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07001_ _01461_ _01921_ _01699_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08952_ rvsingle.dp.rf.rf\[13\]\[25\] _03857_ _01856_ VGND VGND VPWR VPWR _03873_
+ sky130_fd_sc_hd__o21ai_1
X_07903_ _02820_ _02821_ _02822_ _02823_ _01444_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__o221ai_4
X_08883_ _01417_ rvsingle.dp.rf.rf\[16\]\[24\] VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__or2_1
X_07834_ rvsingle.dp.rf.rf\[9\]\[2\] _01539_ _01542_ _02754_ VGND VGND VPWR VPWR _02755_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07765_ _02683_ _01437_ _01721_ _02685_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_79_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06716_ rvsingle.dp.rf.rf\[3\]\[20\] _01255_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09504_ _01962_ _02212_ _03280_ _03255_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07696_ _01096_ rvsingle.dp.rf.rf\[12\]\[5\] _01103_ VGND VGND VPWR VPWR _02617_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09435_ _02848_ _02803_ _02850_ _04142_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__o211a_1
X_06647_ rvsingle.dp.rf.rf\[3\]\[21\] _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__or2b_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ _01185_ _02261_ _02013_ _01959_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06578_ _01498_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__buf_8
XFILLER_0_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08317_ _01878_ rvsingle.dp.rf.rf\[8\]\[8\] VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09297_ _02015_ _02016_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__nand2_1
XANTENNA_40 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_51 ReadData[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_62 ReadData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 ReadData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _01315_ _03161_ _03168_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_84 ReadData[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_95 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08179_ rvsingle.dp.rf.rf\[13\]\[11\] _02379_ _01542_ VGND VGND VPWR VPWR _03100_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_133_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10210_ _04972_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__clkbuf_8
X_11190_ _05377_ net740 _05528_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__mux2_1
X_10141_ _04755_ rvsingle.dp.rf.rf\[28\]\[3\] _04930_ VGND VGND VPWR VPWR _04933_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10072_ _02908_ DataAdr[26] _04872_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10974_ _05314_ _05415_ _05416_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12713_ clknet_leaf_127_clk _00171_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12644_ clknet_leaf_107_clk _00102_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12575_ clknet_leaf_2_clk _00033_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11526_ _04897_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__buf_2
XFILLER_0_108_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11457_ _05639_ net380 _05668_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10408_ _05007_ _05085_ _05065_ net130 VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_22_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11388_ _05640_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ clknet_leaf_92_clk _00585_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10339_ _04859_ net320 _05044_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__mux2_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ clknet_leaf_129_clk _00516_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_12009_ net29 VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07550_ _01592_ _02402_ _02426_ _01481_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__nand4_1
XFILLER_0_49_807 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06501_ _01206_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__buf_8
X_07481_ _02389_ _02401_ _01146_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__nand3_4
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09220_ _04130_ _04132_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__nand3_4
XFILLER_0_158_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06432_ _01352_ _01353_ _01231_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09151_ rvsingle.dp.rf.rf\[2\]\[31\] rvsingle.dp.rf.rf\[3\]\[31\] _01196_ VGND VGND
+ VPWR VPWR _04071_ sky130_fd_sc_hd__mux2_1
X_06363_ _01134_ _01281_ _01283_ _01285_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08102_ _01769_ rvsingle.dp.rf.rf\[22\]\[1\] _01604_ _03022_ VGND VGND VPWR VPWR
+ _03023_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09082_ _01223_ _03988_ _03992_ _01317_ _04001_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__o311a_2
XFILLER_0_44_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06294_ _01216_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__buf_6
XFILLER_0_31_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08033_ _01423_ rvsingle.dp.rf.rf\[3\]\[0\] _01427_ _02953_ VGND VGND VPWR VPWR _02954_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold800 rvsingle.dp.rf.rf\[29\]\[25\] VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 rvsingle.dp.rf.rf\[23\]\[21\] VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09984_ _04713_ _04245_ _04268_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08935_ _01127_ rvsingle.dp.rf.rf\[2\]\[25\] VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08866_ rvsingle.dp.rf.rf\[30\]\[24\] rvsingle.dp.rf.rf\[31\]\[24\] _01658_ VGND
+ VGND VPWR VPWR _03787_ sky130_fd_sc_hd__mux2_1
X_07817_ _02736_ _02737_ _01502_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__o21ai_1
X_08797_ _03715_ _01689_ _02273_ _03717_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__a211o_1
XFILLER_0_169_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07748_ rvsingle.dp.rf.rf\[0\]\[3\] rvsingle.dp.rf.rf\[1\]\[3\] _01241_ VGND VGND
+ VPWR VPWR _02669_ sky130_fd_sc_hd__mux2_1
X_07679_ rvsingle.dp.rf.rf\[20\]\[5\] rvsingle.dp.rf.rf\[21\]\[5\] rvsingle.dp.rf.rf\[22\]\[5\]
+ rvsingle.dp.rf.rf\[23\]\[5\] _02450_ _01455_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09418_ _03398_ _03402_ _04247_ _03366_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__a211o_1
X_10690_ _05248_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09349_ _01248_ _03467_ _03481_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12360_ net25 VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11311_ _05598_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12291_ _04908_ _04912_ _06070_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__o21ai_1
X_11242_ _05560_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11173_ _05187_ net361 _05511_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10124_ Instr[8] VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10055_ _04858_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__buf_2
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10957_ _05406_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10888_ _04908_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__buf_2
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12627_ clknet_leaf_35_clk _00085_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12558_ clknet_leaf_68_clk _01042_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11509_ _05400_ net569 _05706_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12489_ clknet_leaf_96_clk _00973_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold107 rvsingle.dp.rf.rf\[19\]\[9\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 rvsingle.dp.rf.rf\[1\]\[3\] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 rvsingle.dp.rf.rf\[5\]\[6\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ rvsingle.dp.rf.rf\[19\]\[22\] _01901_ _01244_ VGND VGND VPWR VPWR _01902_
+ sky130_fd_sc_hd__o21ai_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _01660_ _03637_ _03638_ _02410_ _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__o311ai_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _03568_ _03569_ _03454_ _03571_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__o22ai_4
X_07602_ rvsingle.dp.rf.rf\[25\]\[4\] _01602_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08582_ _01422_ _03502_ _01221_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07533_ _01207_ _02453_ _02438_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07464_ rvsingle.dp.rf.rf\[31\]\[6\] _01613_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06415_ _01336_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__buf_4
XFILLER_0_63_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09203_ _01059_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07395_ _02301_ _02314_ _02315_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__nand3_1
XFILLER_0_162_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09134_ _04002_ _04013_ _04051_ _04052_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06346_ _01268_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__buf_4
XFILLER_0_72_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09065_ rvsingle.dp.rf.rf\[3\]\[26\] _01297_ _01302_ VGND VGND VPWR VPWR _03985_
+ sky130_fd_sc_hd__o21a_1
X_06277_ _01199_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__buf_6
XFILLER_0_170_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08016_ _02934_ _01172_ _02936_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__nand3_1
XFILLER_0_102_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold630 rvsingle.dp.rf.rf\[21\]\[17\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold641 rvsingle.dp.rf.rf\[1\]\[28\] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 rvsingle.dp.rf.rf\[17\]\[29\] VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 rvsingle.dp.rf.rf\[12\]\[12\] VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 rvsingle.dp.rf.rf\[0\]\[20\] VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 rvsingle.dp.rf.rf\[20\]\[19\] VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold696 rvsingle.dp.rf.rf\[23\]\[12\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ DataAdr[10] ReadData[10] _04750_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__mux2_1
X_08918_ _01796_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__buf_4
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _04722_ _04723_ _04724_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__nor3_2
XFILLER_0_85_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08849_ _01453_ _01480_ _01579_ _01582_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__o22a_1
XFILLER_0_169_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _05713_ net784 _05885_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__mux2_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _05314_ _05315_ _05317_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__a21oi_1
X_11791_ _05854_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10742_ _05277_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10673_ _05239_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12412_ clknet_leaf_147_clk _00896_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13392_ clknet_leaf_55_clk _00820_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12343_ _06123_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12274_ _06074_ net96 _05178_ _05832_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11225_ _05551_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11156_ _05400_ net793 _05511_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10107_ _04903_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__clkbuf_4
X_11087_ _05398_ rvsingle.dp.rf.rf\[17\]\[20\] _05469_ VGND VGND VPWR VPWR _05478_
+ sky130_fd_sc_hd__mux2_1
X_10038_ _01169_ _02259_ _01170_ _04599_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__or4_2
XFILLER_0_72_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11989_ net182 _05940_ _05835_ _05513_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_129_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06200_ Instr[20] VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07180_ _02015_ _02016_ _02098_ _02100_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__and4_2
XFILLER_0_171_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09821_ _04650_ _04653_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09752_ _04590_ PC[20] VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__and2_1
X_06964_ _01098_ rvsingle.dp.rf.rf\[18\]\[22\] VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__nor2_1
X_08703_ _01499_ rvsingle.dp.rf.rf\[8\]\[14\] _03623_ _01496_ VGND VGND VPWR VPWR
+ _03624_ sky130_fd_sc_hd__o211ai_1
X_06895_ _01336_ rvsingle.dp.rf.rf\[6\]\[23\] VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__nor2_1
X_09683_ _04509_ _04517_ _04516_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08634_ _01545_ rvsingle.dp.rf.rf\[24\]\[12\] _02395_ VGND VGND VPWR VPWR _03555_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _02303_ rvsingle.dp.rf.rf\[3\]\[12\] _01953_ _03485_ VGND VGND VPWR VPWR
+ _03486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07516_ rvsingle.dp.rf.rf\[12\]\[6\] rvsingle.dp.rf.rf\[13\]\[6\] rvsingle.dp.rf.rf\[14\]\[6\]
+ rvsingle.dp.rf.rf\[15\]\[6\] _01462_ _01727_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__mux4_2
X_08496_ _03408_ _03411_ _02491_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07447_ _02117_ rvsingle.dp.rf.rf\[18\]\[7\] _01654_ _02367_ VGND VGND VPWR VPWR
+ _02368_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07378_ _02297_ _01691_ _01727_ _02298_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06329_ rvsingle.dp.rf.rf\[1\]\[29\] _01089_ _01093_ _01251_ VGND VGND VPWR VPWR
+ _01252_ sky130_fd_sc_hd__o211ai_1
X_09117_ _01127_ rvsingle.dp.rf.rf\[16\]\[26\] VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09048_ _03857_ rvsingle.dp.rf.rf\[11\]\[27\] _03967_ VGND VGND VPWR VPWR _03968_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold460 rvsingle.dp.rf.rf\[16\]\[23\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 rvsingle.dp.rf.rf\[17\]\[1\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _05291_ rvsingle.dp.rf.rf\[31\]\[16\] _05431_ VGND VGND VPWR VPWR _05437_
+ sky130_fd_sc_hd__mux2_1
Xhold482 rvsingle.dp.rf.rf\[0\]\[25\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 rvsingle.dp.rf.rf\[10\]\[13\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ clknet_leaf_140_clk _00419_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _05476_ net543 _05913_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__mux2_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ clknet_leaf_148_clk _00350_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_300 _01603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _04833_ net536 _05874_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__mux2_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11774_ _05837_ net209 _05751_ _05841_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__a22o_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10725_ _05266_ net773 _05257_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__mux2_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10656_ _05187_ net402 _05219_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13375_ clknet_leaf_133_clk _00803_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10587_ _05189_ _05143_ _05190_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12326_ _06114_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12257_ _05744_ net231 _06074_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11208_ _05207_ net534 _05541_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__mux2_1
X_12188_ _06060_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
X_11139_ _05209_ rvsingle.dp.rf.rf\[16\]\[13\] _05499_ VGND VGND VPWR VPWR _05505_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06680_ _01597_ _01598_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08350_ rvsingle.dp.rf.rf\[19\]\[8\] _01877_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07301_ _02219_ _02221_ _01512_ _01116_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08281_ _01618_ rvsingle.dp.rf.rf\[20\]\[10\] _01489_ VGND VGND VPWR VPWR _03202_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07232_ _01482_ _01171_ _01584_ _02152_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_128_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07163_ rvsingle.dp.rf.rf\[21\]\[18\] _01296_ _01309_ VGND VGND VPWR VPWR _02084_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07094_ _01959_ _02012_ _02014_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__nand3_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ PC[23] PC[24] _04612_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__and3_1
X_07996_ rvsingle.dp.rf.rf\[27\]\[0\] _01240_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__and2b_1
X_09735_ _04454_ _04455_ _04575_ _04459_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__o211ai_1
X_06947_ _01864_ _01867_ _01112_ _01116_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09666_ PC[12] _04500_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__xor2_2
X_06878_ _01796_ rvsingle.dp.rf.rf\[21\]\[23\] _01798_ VGND VGND VPWR VPWR _01799_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _01878_ rvsingle.dp.rf.rf\[20\]\[12\] VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__nor2_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09597_ _04447_ _04448_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__nand2_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ rvsingle.dp.rf.rf\[12\]\[13\] rvsingle.dp.rf.rf\[13\]\[13\] _01468_ VGND
+ VGND VPWR VPWR _03469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_143_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_143_clk sky130_fd_sc_hd__clkbuf_16
X_08479_ _02505_ _03341_ _03364_ _02375_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10510_ _05144_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11490_ _04795_ net663 _05695_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10441_ _05105_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_985 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13160_ clknet_leaf_103_clk _00618_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10372_ _05058_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__buf_8
XFILLER_0_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12111_ _06025_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13091_ clknet_leaf_120_clk _00549_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_12042_ _04807_ net530 _05983_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__mux2_1
Xhold290 rvsingle.dp.rf.rf\[17\]\[17\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ clknet_leaf_51_clk _00402_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12875_ clknet_leaf_88_clk _00333_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _01567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 _01620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_163 _01695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11826_ _05862_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__buf_6
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_185 _01901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 _03644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11757_ _05842_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_134_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_134_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10708_ _04846_ rvsingle.dp.rf.rf\[21\]\[21\] _05257_ VGND VGND VPWR VPWR _05258_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11688_ _05740_ net632 _05795_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10639_ _05220_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13358_ clknet_leaf_68_clk _00786_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12309_ _06105_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__clkbuf_1
X_13289_ clknet_leaf_99_clk _00747_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07850_ _01148_ rvsingle.dp.rf.rf\[6\]\[2\] _01611_ _02770_ VGND VGND VPWR VPWR _02771_
+ sky130_fd_sc_hd__o211ai_1
X_06801_ _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07781_ _01087_ rvsingle.dp.rf.rf\[11\]\[3\] _01611_ _02701_ VGND VGND VPWR VPWR
+ _02702_ sky130_fd_sc_hd__o211ai_1
X_09520_ _04340_ _04395_ VGND VGND VPWR VPWR DataAdr[1] sky130_fd_sc_hd__nand2_8
X_06732_ _01644_ _01649_ _01652_ _01503_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06663_ _01183_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__buf_4
X_09451_ _04310_ _04356_ _04136_ _04357_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_94_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08402_ _01562_ rvsingle.dp.rf.rf\[10\]\[9\] _01620_ _03322_ VGND VGND VPWR VPWR
+ _03323_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06594_ rvsingle.dp.rf.rf\[29\]\[21\] _01488_ _01497_ _01514_ VGND VGND VPWR VPWR
+ _01515_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_59_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09382_ _03227_ _03221_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08333_ _01853_ _03248_ _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_125_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_125_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_145_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08264_ _03183_ _03184_ _02351_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07215_ _02132_ _02133_ _01503_ _02135_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__o211ai_2
X_08195_ _02302_ _03115_ _01699_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_116_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07146_ _02064_ _01870_ _01153_ _02041_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__nand4_1
XFILLER_0_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07077_ _01614_ rvsingle.dp.rf.rf\[0\]\[19\] VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07979_ _02896_ _02897_ _02898_ _02899_ _01600_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09718_ _04558_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__or2b_1
X_10990_ _05381_ net355 _05419_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09649_ _04481_ _04489_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a21oi_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12660_ clknet_leaf_59_clk _00118_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _04904_ _05766_ _05146_ _05767_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_116_clk sky130_fd_sc_hd__clkbuf_16
X_12591_ clknet_leaf_37_clk _00049_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11542_ _05727_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11473_ _05377_ net623 _05684_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__mux2_1
X_13212_ clknet_leaf_14_clk _00670_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10424_ _05093_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_9_clk _00601_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10355_ net84 VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _04909_ _04913_ _04969_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__o21ai_1
X_13074_ clknet_leaf_57_clk _00532_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12025_ _04764_ net585 _05976_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12927_ clknet_leaf_2_clk _00385_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12858_ clknet_leaf_4_clk _00316_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11809_ _05865_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_107_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_107_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12789_ clknet_leaf_64_clk _00247_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07000_ rvsingle.dp.rf.rf\[4\]\[22\] rvsingle.dp.rf.rf\[5\]\[22\] rvsingle.dp.rf.rf\[6\]\[22\]
+ rvsingle.dp.rf.rf\[7\]\[22\] _01335_ _01199_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08951_ _01257_ rvsingle.dp.rf.rf\[12\]\[25\] VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07902_ rvsingle.dp.rf.rf\[5\]\[2\] _01687_ _02268_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__o21ai_1
X_08882_ _01179_ _03802_ _01184_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07833_ _01381_ rvsingle.dp.rf.rf\[8\]\[2\] VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__or2_1
X_07764_ _01827_ rvsingle.dp.rf.rf\[23\]\[3\] _01808_ _02684_ VGND VGND VPWR VPWR
+ _02685_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09503_ _04388_ VGND VGND VPWR VPWR WriteData[9] sky130_fd_sc_hd__clkbuf_4
X_06715_ rvsingle.dp.rf.rf\[1\]\[20\] _01148_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07695_ rvsingle.dp.rf.rf\[15\]\[5\] _01779_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__and2b_1
X_09434_ _04151_ _04334_ _04125_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__a21oi_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06646_ _01566_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__buf_8
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09365_ _04214_ _04280_ _04213_ _02100_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06577_ Instr[20] VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__buf_6
XFILLER_0_118_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08316_ _03233_ _03234_ _03235_ _03236_ _02488_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_47_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09296_ _01737_ _01740_ _04143_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__o21ai_2
XANTENNA_30 Instr[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 ReadData[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 ReadData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08247_ _01422_ _03162_ _03167_ _01699_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__o211ai_1
XANTENNA_74 ReadData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 ReadData[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08178_ _01545_ rvsingle.dp.rf.rf\[12\]\[11\] VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07129_ _01559_ rvsingle.dp.rf.rf\[0\]\[18\] _02049_ _01543_ VGND VGND VPWR VPWR
+ _02050_ sky130_fd_sc_hd__o211ai_1
X_10140_ _04932_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10071_ _02909_ _02799_ _02910_ ReadData[26] _04245_ VGND VGND VPWR VPWR _04872_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_159_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10973_ net112 _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12712_ clknet_leaf_104_clk _00170_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12643_ clknet_leaf_115_clk _00101_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12574_ clknet_leaf_146_clk _00032_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11525_ _05715_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11456_ _05677_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10407_ _05006_ _05068_ _05069_ _05065_ net6 VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__a32o_1
XFILLER_0_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11387_ _05639_ net295 _05629_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13126_ clknet_leaf_111_clk _00584_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _05046_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__clkbuf_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ clknet_leaf_126_clk _00515_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10269_ _04859_ net322 _05001_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12008_ _05970_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06500_ rvsingle.dp.rf.rf\[28\]\[21\] rvsingle.dp.rf.rf\[29\]\[21\] _01420_ VGND
+ VGND VPWR VPWR _01421_ sky130_fd_sc_hd__mux2_1
X_07480_ _01156_ _02394_ _02400_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__nand3_1
XFILLER_0_159_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06431_ rvsingle.dp.rf.rf\[20\]\[28\] rvsingle.dp.rf.rf\[21\]\[28\] rvsingle.dp.rf.rf\[22\]\[28\]
+ rvsingle.dp.rf.rf\[23\]\[28\] _01338_ _01303_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06362_ _01133_ _01284_ _01117_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09150_ rvsingle.dp.rf.rf\[4\]\[31\] rvsingle.dp.rf.rf\[5\]\[31\] rvsingle.dp.rf.rf\[6\]\[31\]
+ rvsingle.dp.rf.rf\[7\]\[31\] _01225_ _01203_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_671 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08101_ rvsingle.dp.rf.rf\[23\]\[1\] _01124_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__or2b_1
XFILLER_0_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09081_ _02191_ _03994_ _03996_ _01219_ _04000_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__a311o_1
XFILLER_0_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06293_ _01215_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__inv_4
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08032_ _01425_ rvsingle.dp.rf.rf\[2\]\[0\] VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold801 rvsingle.dp.rf.rf\[13\]\[20\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold812 rvsingle.dp.rf.rf\[31\]\[15\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09983_ _04797_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
X_08934_ _03843_ _03854_ _01147_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08865_ rvsingle.dp.rf.rf\[29\]\[24\] _01540_ _01543_ _03785_ VGND VGND VPWR VPWR
+ _03786_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07816_ rvsingle.dp.rf.rf\[21\]\[3\] _02627_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__and2b_1
X_08796_ _02929_ rvsingle.dp.rf.rf\[11\]\[15\] _01727_ _03716_ VGND VGND VPWR VPWR
+ _03717_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07747_ _02476_ _02577_ _02661_ _02667_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__nand4_2
XFILLER_0_95_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07678_ _02302_ _02594_ _02438_ _02598_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__o211ai_1
X_09417_ _03313_ _04326_ _04325_ _04125_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__a31o_1
X_06629_ rvsingle.dp.rf.rf\[9\]\[21\] _01540_ _01543_ VGND VGND VPWR VPWR _01550_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09348_ _04222_ _04263_ _04257_ _04261_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09279_ _03984_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11310_ _05307_ rvsingle.dp.rf.rf\[15\]\[27\] _05591_ VGND VGND VPWR VPWR _05598_
+ sky130_fd_sc_hd__mux2_1
X_12290_ net90 VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11241_ _05359_ net291 _05552_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11172_ _05521_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__clkbuf_1
X_10123_ _04917_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__buf_2
X_10054_ _04426_ _04616_ _04857_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10956_ _05304_ net510 _05401_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10887_ net73 VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__inv_2
X_12626_ clknet_leaf_41_clk _00084_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12557_ clknet_leaf_43_clk _01041_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11508_ _05683_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__buf_6
XFILLER_0_124_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12488_ clknet_leaf_106_clk _00972_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold108 rvsingle.dp.rf.rf\[17\]\[0\] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold119 rvsingle.dp.rf.rf\[7\]\[22\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ _05400_ rvsingle.dp.rf.rf\[13\]\[21\] _05668_ VGND VGND VPWR VPWR _05669_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ clknet_leaf_65_clk _00567_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _01294_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__buf_6
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08650_ _01960_ _02102_ _02261_ _03570_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__a2bb2oi_1
X_07601_ _02030_ rvsingle.dp.rf.rf\[24\]\[4\] VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08581_ rvsingle.dp.rf.rf\[28\]\[12\] rvsingle.dp.rf.rf\[29\]\[12\] rvsingle.dp.rf.rf\[30\]\[12\]
+ rvsingle.dp.rf.rf\[31\]\[12\] _01416_ _01300_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07532_ rvsingle.dp.rf.rf\[28\]\[6\] rvsingle.dp.rf.rf\[29\]\[6\] rvsingle.dp.rf.rf\[30\]\[6\]
+ rvsingle.dp.rf.rf\[31\]\[6\] _01462_ _01470_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07463_ _02117_ rvsingle.dp.rf.rf\[30\]\[6\] VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09202_ _01063_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__clkbuf_4
X_06414_ _01335_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07394_ Instr[19] VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__buf_8
XFILLER_0_60_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09133_ _04002_ _04013_ _04051_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__nor4_4
XFILLER_0_146_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06345_ _01267_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06276_ _01198_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__buf_6
X_09064_ _03982_ _03983_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__or2b_2
XFILLER_0_142_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08015_ rvsingle.dp.rf.rf\[23\]\[0\] _02929_ _02935_ VGND VGND VPWR VPWR _02936_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold620 rvsingle.dp.rf.rf\[5\]\[25\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold631 rvsingle.dp.rf.rf\[12\]\[25\] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 rvsingle.dp.rf.rf\[0\]\[18\] VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold653 rvsingle.dp.rf.rf\[12\]\[10\] VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 rvsingle.dp.rf.rf\[9\]\[16\] VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 rvsingle.dp.rf.rf\[23\]\[15\] VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 rvsingle.dp.rf.rf\[12\]\[8\] VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold697 rvsingle.dp.rf.rf\[13\]\[14\] VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _04783_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
X_08917_ _01257_ rvsingle.dp.rf.rf\[30\]\[25\] VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__nor2_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ Instr[9] VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__clkbuf_4
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08848_ _01931_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__nand2_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ rvsingle.dp.rf.rf\[24\]\[15\] rvsingle.dp.rf.rf\[25\]\[15\] rvsingle.dp.rf.rf\[26\]\[15\]
+ rvsingle.dp.rf.rf\[27\]\[15\] _01691_ _01244_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__mux4_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _05316_ _05145_ net4 VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__a21oi_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _05713_ net497 _05845_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__mux2_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10741_ _04755_ rvsingle.dp.rf.rf\[20\]\[3\] _05274_ VGND VGND VPWR VPWR _05277_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10672_ _04760_ rvsingle.dp.rf.rf\[21\]\[4\] _05235_ VGND VGND VPWR VPWR _05239_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12411_ clknet_leaf_142_clk _00895_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13391_ clknet_leaf_39_clk _00819_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12342_ _04852_ net574 _06121_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12273_ _05177_ _05835_ _06077_ net171 VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__a2bb2o_1
X_11224_ _05398_ net705 _05541_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11155_ _05490_ net16 _05371_ _05513_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__o2bb2ai_1
X_10106_ _04365_ _04901_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__o21ai_2
X_11086_ _05175_ _05471_ _05463_ net137 VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_87_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
X_10037_ _02908_ DataAdr[21] _04842_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11988_ _05961_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10939_ _04828_ net614 _05387_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12609_ clknet_leaf_140_clk _00067_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09820_ _04651_ _04652_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__nand2_1
X_09751_ Instr[31] VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__buf_2
X_06963_ _01883_ _01526_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_78_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
X_08702_ rvsingle.dp.rf.rf\[9\]\[14\] _01498_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09682_ _04494_ _04497_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__o21bai_2
X_06894_ rvsingle.dp.rf.rf\[5\]\[23\] _01688_ _01689_ VGND VGND VPWR VPWR _01815_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08633_ rvsingle.dp.rf.rf\[25\]\[12\] _01769_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _01468_ rvsingle.dp.rf.rf\[2\]\[12\] VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07515_ _02433_ _01689_ _01702_ _02435_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__a211oi_2
X_08495_ _03412_ _03413_ _03415_ _02323_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07446_ rvsingle.dp.rf.rf\[19\]\[7\] _01557_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_162_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07377_ _01416_ rvsingle.dp.rf.rf\[24\]\[7\] VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09116_ _04033_ _04035_ _01512_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06328_ _01099_ rvsingle.dp.rf.rf\[0\]\[29\] VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09047_ _01744_ rvsingle.dp.rf.rf\[10\]\[27\] _01105_ VGND VGND VPWR VPWR _03967_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06259_ _01066_ _01075_ _01181_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__or3b_2
XFILLER_0_41_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold450 rvsingle.dp.rf.rf\[0\]\[11\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 rvsingle.dp.rf.rf\[20\]\[29\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 rvsingle.dp.rf.rf\[0\]\[19\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 rvsingle.dp.rf.rf\[19\]\[2\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 rvsingle.dp.rf.rf\[5\]\[18\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
X_09949_ _04769_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12960_ clknet_leaf_115_clk _00418_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _05919_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__clkbuf_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ clknet_leaf_141_clk _00349_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 _01603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _05882_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11773_ _05781_ _05847_ _05840_ net153 VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _04897_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__buf_2
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10655_ _05228_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13374_ clknet_leaf_14_clk _00802_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10586_ _04909_ _04913_ _05143_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12325_ _04807_ net804 _06110_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12256_ _06077_ net52 _05164_ _05832_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11207_ _05542_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12187_ _05132_ net378 _06048_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__mux2_1
X_11138_ _05504_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__clkbuf_1
X_11069_ _05459_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_0_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07300_ _01383_ rvsingle.dp.rf.rf\[22\]\[16\] _01260_ _02220_ VGND VGND VPWR VPWR
+ _02221_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_46_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08280_ rvsingle.dp.rf.rf\[23\]\[10\] _01743_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07231_ _01592_ _02149_ _02126_ _01178_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__a31o_1
XFILLER_0_171_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07162_ _01330_ rvsingle.dp.rf.rf\[20\]\[18\] VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07093_ _01482_ _01171_ _01584_ _02013_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09803_ _04635_ _04637_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07995_ _01903_ rvsingle.dp.rf.rf\[26\]\[0\] VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__nor2_4
X_09734_ PC[18] _04564_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__xnor2_1
X_06946_ rvsingle.dp.rf.rf\[5\]\[22\] _01865_ _01759_ _01866_ VGND VGND VPWR VPWR
+ _01867_ sky130_fd_sc_hd__o211ai_1
X_09665_ _04504_ _04511_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06877_ _01797_ rvsingle.dp.rf.rf\[20\]\[23\] _01604_ VGND VGND VPWR VPWR _01798_
+ sky130_fd_sc_hd__o21ba_1
X_08616_ _01377_ _03524_ _03536_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__nand3_4
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ Instr[27] PC[7] VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08547_ rvsingle.dp.rf.rf\[8\]\[13\] rvsingle.dp.rf.rf\[9\]\[13\] rvsingle.dp.rf.rf\[10\]\[13\]
+ rvsingle.dp.rf.rf\[11\]\[13\] _01241_ _01953_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__mux4_2
XFILLER_0_166_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08478_ _03366_ _03367_ _03398_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07429_ rvsingle.dp.rf.rf\[27\]\[7\] _01602_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__and2b_1
XFILLER_0_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10440_ _04747_ rvsingle.dp.rf.rf\[24\]\[2\] _05103_ VGND VGND VPWR VPWR _05105_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10371_ _05067_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12110_ _04807_ net531 _06019_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13090_ clknet_leaf_129_clk _00548_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12041_ _05988_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__clkbuf_1
Xhold280 rvsingle.dp.rf.rf\[1\]\[1\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold291 rvsingle.dp.rf.rf\[29\]\[28\] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ clknet_leaf_40_clk _00401_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _01452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12874_ clknet_leaf_81_clk _00332_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _01567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_153 _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11825_ _05873_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_164 _01695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _01763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_186 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_197 _04210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _05534_ rvsingle.dp.rf.rf\[7\]\[5\] _05837_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10707_ _05234_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__buf_8
XFILLER_0_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11687_ _05802_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10638_ _04846_ net347 _05219_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13357_ clknet_leaf_45_clk _00785_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10569_ _04863_ net254 _05151_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12308_ _04769_ net749 _06099_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__mux2_1
X_13288_ clknet_leaf_121_clk _00746_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12239_ _06072_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__buf_8
XFILLER_0_78_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06800_ _01206_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__buf_6
X_07780_ _01752_ rvsingle.dp.rf.rf\[10\]\[3\] VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06731_ rvsingle.dp.rf.rf\[29\]\[20\] _01646_ _01092_ _01651_ VGND VGND VPWR VPWR
+ _01652_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09450_ _02463_ _02472_ _02432_ _04142_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__o211a_1
X_06662_ _01453_ _01480_ _01579_ _01582_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08401_ rvsingle.dp.rf.rf\[11\]\[9\] _03258_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__or2b_1
XFILLER_0_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09381_ _03064_ _04295_ _03399_ _03405_ _03749_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__a41o_1
X_06593_ _01513_ rvsingle.dp.rf.rf\[28\]\[21\] VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08332_ _03249_ _03250_ _02488_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08263_ rvsingle.dp.rf.rf\[1\]\[10\] _01743_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07214_ rvsingle.dp.rf.rf\[13\]\[17\] _01865_ _01668_ _02134_ VGND VGND VPWR VPWR
+ _02135_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08194_ rvsingle.dp.rf.rf\[0\]\[11\] rvsingle.dp.rf.rf\[1\]\[11\] rvsingle.dp.rf.rf\[2\]\[11\]
+ rvsingle.dp.rf.rf\[3\]\[11\] _02450_ _01708_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07145_ _01960_ _01075_ _01961_ _02065_ _01587_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_42_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07076_ _01993_ _01996_ _01116_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_113_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07978_ rvsingle.dp.rf.rf\[19\]\[0\] _01677_ _01531_ VGND VGND VPWR VPWR _02899_
+ sky130_fd_sc_hd__o21ai_1
X_09717_ _01232_ _02912_ _01175_ _01171_ PC[17] VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a311o_1
X_06929_ _01848_ rvsingle.dp.rf.rf\[10\]\[22\] _01612_ _01849_ VGND VGND VPWR VPWR
+ _01850_ sky130_fd_sc_hd__o211ai_1
X_09648_ _04494_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__or2_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ Instr[25] _04429_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__or2_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11610_ _04976_ _05417_ _05149_ net564 VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__o31a_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ clknet_leaf_71_clk _00048_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11541_ _05724_ net715 _05726_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11472_ _05687_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13211_ clknet_leaf_17_clk _00669_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10423_ _04898_ net616 _05082_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13142_ clknet_leaf_31_clk _00600_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10354_ _05054_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13073_ clknet_leaf_48_clk _00531_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ net68 VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__inv_2
X_12024_ _05980_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12926_ clknet_leaf_150_clk _00384_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ clknet_leaf_8_clk _00315_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _05728_ net721 _05863_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ clknet_leaf_60_clk _00246_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11739_ _04915_ _04917_ _04965_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13409_ clknet_leaf_139_clk _00837_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08950_ _03867_ _03868_ _03870_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__o21ai_1
X_07901_ _01707_ rvsingle.dp.rf.rf\[4\]\[2\] VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__nor2_1
X_08881_ _01153_ _03790_ _03801_ _01537_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__and4_1
XFILLER_0_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07832_ rvsingle.dp.rf.rf\[11\]\[2\] _01539_ _02337_ VGND VGND VPWR VPWR _02753_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07763_ _01828_ rvsingle.dp.rf.rf\[22\]\[3\] VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__or2_1
X_09502_ _04377_ _03341_ _03364_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__and3_4
XFILLER_0_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06714_ _01614_ rvsingle.dp.rf.rf\[0\]\[20\] VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__nor2_1
X_07694_ _01125_ rvsingle.dp.rf.rf\[14\]\[5\] VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09433_ _04334_ _04151_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__or2_1
X_06645_ _01095_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__buf_6
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _04165_ _02184_ _02265_ _04279_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__a31oi_1
X_06576_ _01496_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08315_ rvsingle.dp.rf.rf\[13\]\[8\] _01487_ _01496_ VGND VGND VPWR VPWR _03236_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09295_ _03741_ _02261_ _03727_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__a21oi_1
XANTENNA_20 DataAdr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 Instr[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 ReadData[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08246_ _03163_ _03164_ _02543_ _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_64 ReadData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_75 ReadData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_86 ReadData[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 ReadData[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08177_ _03095_ _03097_ _02364_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_132_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07128_ rvsingle.dp.rf.rf\[1\]\[18\] _01558_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07059_ _01842_ rvsingle.dp.rf.rf\[29\]\[19\] _01979_ VGND VGND VPWR VPWR _01980_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10070_ _04871_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10972_ _04967_ _04968_ _04925_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__and3_2
X_12711_ clknet_leaf_98_clk _00169_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12642_ clknet_leaf_128_clk _00100_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12573_ clknet_leaf_133_clk _01057_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11524_ _05359_ net309 _05706_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11455_ _05266_ net503 _05668_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10406_ _05005_ _05085_ _05065_ net146 VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ _04903_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13125_ clknet_leaf_101_clk _00583_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10337_ _04853_ net456 _05044_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ clknet_leaf_116_clk _00514_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10268_ _05008_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__clkbuf_1
X_12007_ _05639_ net243 _05960_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10199_ net41 VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12909_ clknet_leaf_43_clk _00367_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06430_ rvsingle.dp.rf.rf\[16\]\[28\] rvsingle.dp.rf.rf\[17\]\[28\] rvsingle.dp.rf.rf\[18\]\[28\]
+ rvsingle.dp.rf.rf\[19\]\[28\] _01338_ _01303_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__mux4_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06361_ rvsingle.dp.rf.rf\[28\]\[29\] rvsingle.dp.rf.rf\[29\]\[29\] rvsingle.dp.rf.rf\[30\]\[29\]
+ rvsingle.dp.rf.rf\[31\]\[29\] _01138_ _01106_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08100_ rvsingle.dp.rf.rf\[21\]\[1\] _01381_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09080_ _03997_ _01310_ _02191_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__a211oi_1
X_06292_ Instr[18] VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08031_ _02950_ _02951_ _01206_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold802 rvsingle.dp.rf.rf\[22\]\[3\] VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold813 rvsingle.dp.rf.rf\[19\]\[21\] VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09982_ _04796_ net519 _04791_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__mux2_1
X_08933_ _01133_ _03848_ _03853_ _01157_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_110_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08864_ _01780_ rvsingle.dp.rf.rf\[28\]\[24\] VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07815_ _01602_ rvsingle.dp.rf.rf\[20\]\[3\] _01258_ VGND VGND VPWR VPWR _02736_
+ sky130_fd_sc_hd__o21bai_1
X_08795_ _01240_ rvsingle.dp.rf.rf\[10\]\[15\] VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__or2_1
X_07746_ _02664_ _02665_ _02666_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__nand3_2
XFILLER_0_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07677_ _02595_ _02285_ _01206_ _02597_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09416_ _03313_ _04325_ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__a21oi_1
X_06628_ _01383_ rvsingle.dp.rf.rf\[8\]\[21\] VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09347_ _04258_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__inv_2
X_06559_ _01316_ _01467_ _01479_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__and3_2
XFILLER_0_63_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09278_ _04002_ _04013_ _04191_ _04055_ _04193_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__o32ai_1
XFILLER_0_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08229_ _01327_ rvsingle.dp.rf.rf\[26\]\[10\] VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11240_ _05559_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11171_ _05266_ net429 _05511_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__mux2_1
X_10122_ _04723_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10053_ _04505_ _01071_ _01079_ _04855_ _04856_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__a32o_1
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10955_ _05405_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10886_ _04904_ _05183_ _05336_ _05362_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12625_ clknet_leaf_48_clk _00083_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12556_ clknet_leaf_51_clk _01040_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11507_ _05705_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12487_ clknet_leaf_101_clk _00971_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold109 rvsingle.dp.rf.rf\[19\]\[0\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11438_ _05645_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__buf_6
XFILLER_0_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11369_ _05630_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ clknet_leaf_61_clk _00566_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13039_ clknet_leaf_57_clk _00497_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07600_ _02517_ _02518_ _02520_ _01617_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__o211ai_1
X_08580_ _03498_ _01309_ _02302_ _03500_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07531_ _02302_ _02451_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07462_ _02378_ _02380_ _02381_ _02382_ _02351_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_159_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09201_ _02907_ _02963_ _02966_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06413_ _01240_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07393_ _02302_ _02305_ _02307_ _02313_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_85_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09132_ _01581_ _04050_ _01837_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06344_ _01135_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09063_ _03979_ _03981_ _03939_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06275_ _01197_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__buf_6
XFILLER_0_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08014_ _01425_ rvsingle.dp.rf.rf\[22\]\[0\] _01197_ VGND VGND VPWR VPWR _02935_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold610 rvsingle.dp.rf.rf\[30\]\[3\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 rvsingle.dp.rf.rf\[29\]\[27\] VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold632 rvsingle.dp.rf.rf\[10\]\[8\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 rvsingle.dp.rf.rf\[6\]\[9\] VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 rvsingle.dp.rf.rf\[17\]\[2\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold665 rvsingle.dp.rf.rf\[6\]\[20\] VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 rvsingle.dp.rf.rf\[2\]\[8\] VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 rvsingle.dp.rf.rf\[2\]\[17\] VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 rvsingle.dp.rf.rf\[31\]\[28\] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _04782_ net538 _04741_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08916_ rvsingle.dp.rf.rf\[29\]\[25\] _01488_ _01497_ VGND VGND VPWR VPWR _03837_
+ sky130_fd_sc_hd__o21ai_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ Instr[10] VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__clkbuf_4
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _03760_ _03765_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__o21ai_2
X_08778_ _01084_ _01171_ _01584_ _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__o211ai_2
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _02648_ _02649_ _01502_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__o21ai_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _05276_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10671_ _05238_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12410_ clknet_leaf_5_clk _00894_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ clknet_leaf_65_clk _00818_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12341_ _06122_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12272_ _06086_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11223_ _05550_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11154_ _04967_ _04968_ _04976_ _04839_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__or4b_2
XFILLER_0_101_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10105_ PC[29] PC[30] _04681_ _04691_ _04425_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__a311o_1
X_11085_ _05463_ net188 _05174_ _05464_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__a22o_1
X_10036_ _02909_ _02799_ _02910_ ReadData[21] _04715_ VGND VGND VPWR VPWR _04842_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11987_ _04833_ net241 _05960_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10938_ _05395_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10869_ _05352_ net238 _05320_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12608_ clknet_leaf_118_clk _00066_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12539_ clknet_leaf_145_clk _01023_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06962_ _01260_ _01876_ _01879_ _01565_ _01882_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__o311ai_1
X_09750_ _04585_ _04552_ _04588_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__o21ai_2
X_08701_ rvsingle.dp.rf.rf\[11\]\[14\] _01487_ _01523_ VGND VGND VPWR VPWR _03622_
+ sky130_fd_sc_hd__o21ai_1
X_09681_ _04509_ _04510_ _04518_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__or3_1
X_06893_ _01336_ rvsingle.dp.rf.rf\[4\]\[23\] VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08632_ _03550_ _02488_ _03552_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08563_ rvsingle.dp.rf.rf\[0\]\[12\] rvsingle.dp.rf.rf\[1\]\[12\] _01691_ VGND VGND
+ VPWR VPWR _03484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07514_ _01440_ rvsingle.dp.rf.rf\[11\]\[6\] _01696_ _02434_ VGND VGND VPWR VPWR
+ _02435_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08494_ _01860_ rvsingle.dp.rf.rf\[29\]\[13\] _03414_ VGND VGND VPWR VPWR _03415_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07445_ rvsingle.dp.rf.rf\[17\]\[7\] _01136_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__and2b_1
XFILLER_0_146_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07376_ rvsingle.dp.rf.rf\[25\]\[7\] VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09115_ rvsingle.dp.rf.rf\[23\]\[26\] _03839_ _04034_ VGND VGND VPWR VPWR _04035_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06327_ _01182_ _01186_ _01249_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__nand3_4
XFILLER_0_162_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09046_ _03963_ _03965_ _03782_ _01506_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06258_ _01085_ WriteData[30] _01180_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold440 rvsingle.dp.rf.rf\[15\]\[29\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ _01112_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_8
Xhold451 rvsingle.dp.rf.rf\[16\]\[27\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 rvsingle.dp.rf.rf\[24\]\[26\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 rvsingle.dp.rf.rf\[14\]\[2\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 rvsingle.dp.rf.rf\[13\]\[9\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 rvsingle.dp.rf.rf\[14\]\[9\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09948_ _04767_ _04444_ _04426_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__a2bb2o_4
X_09879_ _04618_ PC[31] VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__and2_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _05344_ net360 _05913_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__mux2_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ clknet_leaf_5_clk _00348_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_302 _01603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _05173_ rvsingle.dp.rf.rf\[23\]\[18\] _05874_ VGND VGND VPWR VPWR _05882_
+ sky130_fd_sc_hd__mux2_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11772_ _05749_ _05847_ _05840_ net69 VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _05265_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10654_ _04898_ net624 _05219_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13373_ clknet_leaf_144_clk _00801_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10585_ net64 VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__inv_2
X_12324_ _06113_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12255_ _06080_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__clkbuf_1
X_11206_ _05334_ net796 _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__mux2_1
X_12186_ _06059_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_1
X_11137_ _05207_ rvsingle.dp.rf.rf\[16\]\[12\] _05499_ VGND VGND VPWR VPWR _05504_
+ sky130_fd_sc_hd__mux2_1
X_11068_ _05463_ net167 _05164_ _05464_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__a22o_1
X_10019_ _04827_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__buf_2
XFILLER_0_149_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07230_ _01960_ _02102_ _01961_ _02150_ _01587_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_6_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07161_ rvsingle.dp.rf.rf\[16\]\[18\] rvsingle.dp.rf.rf\[17\]\[18\] rvsingle.dp.rf.rf\[18\]\[18\]
+ rvsingle.dp.rf.rf\[19\]\[18\] _01242_ _01434_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07092_ _02011_ _01084_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09802_ _04632_ _04633_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__a21o_1
X_07994_ _02908_ _01067_ _02913_ _02914_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__a22oi_2
X_06945_ _01148_ rvsingle.dp.rf.rf\[4\]\[22\] VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09733_ _04569_ _04573_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__xnor2_1
X_06876_ _01124_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__clkbuf_8
X_09664_ _04509_ _04510_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08615_ _03527_ _03530_ _01156_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09595_ Instr[27] PC[7] VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__nand2_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08546_ _03457_ _03459_ _03466_ _01187_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08477_ _01351_ _01202_ _03382_ _03397_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_9_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07428_ _01658_ rvsingle.dp.rf.rf\[26\]\[7\] _01259_ VGND VGND VPWR VPWR _02349_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07359_ _01460_ _02277_ _02279_ _01216_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10370_ _04747_ net659 _05065_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09029_ rvsingle.dp.rf.rf\[28\]\[27\] rvsingle.dp.rf.rf\[29\]\[27\] rvsingle.dp.rf.rf\[30\]\[27\]
+ rvsingle.dp.rf.rf\[31\]\[27\] _01559_ _03840_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12040_ _04801_ net677 _05983_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold270 rvsingle.dp.rf.rf\[23\]\[8\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 rvsingle.dp.rf.rf\[10\]\[28\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 rvsingle.dp.rf.rf\[6\]\[28\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ clknet_leaf_52_clk _00400_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12873_ clknet_leaf_95_clk _00331_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _01452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _01567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _04785_ net317 _05863_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__mux2_1
XANTENNA_154 _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _01695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _01763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_198 _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _05840_ net36 _05735_ _05841_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10706_ _05256_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__clkbuf_1
X_11686_ _05381_ rvsingle.dp.rf.rf\[10\]\[7\] _05795_ VGND VGND VPWR VPWR _05802_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10637_ _05193_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__buf_8
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13356_ clknet_leaf_67_clk _00784_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10568_ _05179_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_1
X_12307_ _06104_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10499_ _05101_ _05137_ _05103_ net216 VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__a2bb2o_1
X_13287_ clknet_leaf_89_clk _00745_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12238_ _04919_ _04732_ _05835_ _04737_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__or4b_1
X_12169_ _06054_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06730_ _01650_ rvsingle.dp.rf.rf\[28\]\[20\] VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06661_ _01581_ _01578_ _01486_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__a21oi_2
X_08400_ _03319_ _03320_ _02483_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__o21ai_1
X_09380_ _03313_ _03317_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__and2_1
X_06592_ _01267_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__buf_6
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08331_ rvsingle.dp.rf.rf\[5\]\[8\] _02481_ _01496_ _03251_ VGND VGND VPWR VPWR _03252_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_129_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08262_ _01763_ rvsingle.dp.rf.rf\[0\]\[10\] _01604_ VGND VGND VPWR VPWR _03183_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07213_ _01753_ rvsingle.dp.rf.rf\[12\]\[17\] VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08193_ _02093_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07144_ _01962_ _01100_ _02041_ _02064_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07075_ _01994_ _01995_ _01632_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07977_ rvsingle.dp.rf.rf\[18\]\[0\] _01126_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__nor2_1
X_09716_ _04507_ _01176_ PC[17] VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__o21a_1
X_06928_ rvsingle.dp.rf.rf\[11\]\[22\] _01097_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09647_ PC[11] _04493_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__nor2_1
X_06859_ _01779_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__buf_8
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _04430_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08529_ _01520_ _03446_ _03447_ _01502_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11540_ _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__buf_8
XFILLER_0_92_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11471_ _05531_ rvsingle.dp.rf.rf\[12\]\[3\] _05684_ VGND VGND VPWR VPWR _05687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10422_ _05092_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__clkbuf_1
X_13210_ clknet_leaf_21_clk _00668_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10353_ _04904_ net337 _05044_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__mux2_1
X_13141_ clknet_leaf_37_clk _00599_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13072_ clknet_leaf_51_clk _00530_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10284_ _05016_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12023_ _04759_ net396 _05976_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__mux2_1
X_12925_ clknet_leaf_142_clk _00383_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ clknet_leaf_33_clk _00314_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _05864_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ clknet_leaf_27_clk _00245_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11738_ _05828_ _05792_ _05829_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11669_ _04720_ _04728_ _05142_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__and3_2
XFILLER_0_153_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13408_ clknet_leaf_119_clk _00836_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13339_ clknet_leaf_77_clk rvsingle.dp.PCNext\[16\] _00016_ VGND VGND VPWR VPWR PC[16]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07900_ rvsingle.dp.rf.rf\[7\]\[2\] _01687_ _01470_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08880_ _03792_ _03794_ _01378_ _03800_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__o211ai_2
X_07831_ _02030_ rvsingle.dp.rf.rf\[10\]\[2\] VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07762_ rvsingle.dp.rf.rf\[20\]\[3\] rvsingle.dp.rf.rf\[21\]\[3\] _01335_ VGND VGND
+ VPWR VPWR _02683_ sky130_fd_sc_hd__mux2_1
X_09501_ _04387_ VGND VGND VPWR VPWR WriteData[10] sky130_fd_sc_hd__clkbuf_4
X_06713_ _01155_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__clkbuf_8
X_07693_ _02610_ _02611_ _02613_ _02329_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06644_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__clkbuf_8
X_09432_ _04120_ _04338_ _04125_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__a211o_2
XFILLER_0_149_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09363_ _03765_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__inv_2
X_06575_ _01091_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__buf_6
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08314_ _01493_ rvsingle.dp.rf.rf\[12\]\[8\] VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09294_ _01898_ _04123_ _04208_ _04209_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__o31a_4
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_10 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_21 Instr[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_32 Instr[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_43 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08245_ rvsingle.dp.rf.rf\[1\]\[10\] _01295_ _01308_ _03165_ VGND VGND VPWR VPWR
+ _03166_ sky130_fd_sc_hd__o211ai_1
XANTENNA_54 ReadData[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 ReadData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_76 ReadData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_87 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ _01558_ rvsingle.dp.rf.rf\[2\]\[11\] _01880_ _03096_ VGND VGND VPWR VPWR
+ _03097_ sky130_fd_sc_hd__o211a_1
XANTENNA_98 ReadData[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07127_ _01559_ rvsingle.dp.rf.rf\[2\]\[18\] _01260_ _02047_ VGND VGND VPWR VPWR
+ _02048_ sky130_fd_sc_hd__o211ai_1
X_07058_ _01675_ rvsingle.dp.rf.rf\[28\]\[19\] _01104_ VGND VGND VPWR VPWR _01979_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10971_ _05413_ _05368_ _05414_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12710_ clknet_leaf_115_clk _00168_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12641_ clknet_leaf_140_clk _00099_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12572_ clknet_leaf_150_clk _01056_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11523_ _05714_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11454_ _05676_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_807 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10405_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__clkbuf_8
X_11385_ _05638_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13124_ clknet_leaf_124_clk _00582_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10336_ _05045_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__clkbuf_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _04853_ rvsingle.dp.rf.rf\[27\]\[22\] _05001_ VGND VGND VPWR VPWR _05008_
+ sky130_fd_sc_hd__mux2_1
X_13055_ clknet_leaf_13_clk _00513_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_12006_ _05969_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10198_ _04962_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12908_ clknet_leaf_50_clk _00366_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12839_ clknet_leaf_98_clk _00297_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06360_ rvsingle.dp.rf.rf\[25\]\[29\] _01090_ _01094_ _01282_ VGND VGND VPWR VPWR
+ _01283_ sky130_fd_sc_hd__o211ai_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06291_ _01212_ _01213_ _01210_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08030_ rvsingle.dp.rf.rf\[1\]\[0\] _01690_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold803 rvsingle.dp.rf.rf\[15\]\[16\] VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold814 rvsingle.dp.rf.rf\[8\]\[27\] VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09981_ _04795_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08932_ _03849_ _03850_ _03852_ _02236_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__o211ai_1
X_08863_ rvsingle.dp.rf.rf\[24\]\[24\] rvsingle.dp.rf.rf\[25\]\[24\] rvsingle.dp.rf.rf\[26\]\[24\]
+ rvsingle.dp.rf.rf\[27\]\[24\] _01137_ _01612_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__mux4_2
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07814_ _02733_ _02030_ _01542_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__a211oi_1
X_08794_ rvsingle.dp.rf.rf\[8\]\[15\] rvsingle.dp.rf.rf\[9\]\[15\] _02440_ VGND VGND
+ VPWR VPWR _03715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07745_ _01065_ _01074_ _01178_ _02662_ _02609_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_74_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07676_ _01294_ rvsingle.dp.rf.rf\[31\]\[5\] _01243_ _02596_ VGND VGND VPWR VPWR
+ _02597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09415_ _03399_ _03405_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__nand2_1
X_06627_ _01538_ _01541_ _01547_ _01512_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_164_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06558_ _01230_ _01472_ _01474_ _01477_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__o221ai_1
X_09346_ _04257_ _04260_ _04261_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09277_ _03908_ _04192_ _03775_ _03910_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__a22oi_4
X_06489_ _01347_ _01288_ _01290_ _01409_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08228_ rvsingle.dp.rf.rf\[24\]\[10\] rvsingle.dp.rf.rf\[25\]\[10\] _01349_ VGND
+ VGND VPWR VPWR _03149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08159_ _01630_ rvsingle.dp.rf.rf\[26\]\[11\] _01259_ _03079_ VGND VGND VPWR VPWR
+ _03080_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11170_ _05520_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10121_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__clkbuf_2
X_10052_ _02908_ DataAdr[23] VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10954_ _05354_ net781 _05401_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10885_ _05337_ _05338_ _05339_ _05084_ net300 VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__o41a_1
XFILLER_0_156_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12624_ clknet_leaf_70_clk _00082_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12555_ clknet_leaf_88_clk _01039_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11506_ _05398_ net736 _05695_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12486_ clknet_leaf_108_clk _00970_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11437_ _05667_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11368_ _05400_ net810 _05629_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ clknet_leaf_16_clk _00565_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _05036_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__clkbuf_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _05592_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__clkbuf_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ clknet_4_15_0_clk _00496_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07530_ rvsingle.dp.rf.rf\[24\]\[6\] rvsingle.dp.rf.rf\[25\]\[6\] rvsingle.dp.rf.rf\[26\]\[6\]
+ rvsingle.dp.rf.rf\[27\]\[6\] _02450_ _01455_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07461_ rvsingle.dp.rf.rf\[25\]\[6\] _01539_ _01542_ VGND VGND VPWR VPWR _02382_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06412_ _01231_ _01325_ _01333_ _01223_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__o211a_1
X_09200_ _01250_ _04063_ _04114_ _04115_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__o2bb2ai_4
X_07392_ _02310_ _02312_ _02291_ _01446_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06343_ rvsingle.dp.rf.rf\[13\]\[29\] _01089_ _01093_ _01265_ VGND VGND VPWR VPWR
+ _01266_ sky130_fd_sc_hd__o211a_1
X_09131_ _01066_ _01075_ _01482_ _01483_ _04050_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__o221a_2
XFILLER_0_72_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09062_ _03939_ _03979_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nor3_2
X_06274_ Instr[16] VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__buf_4
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08013_ rvsingle.dp.rf.rf\[21\]\[0\] _02929_ _01307_ _02933_ VGND VGND VPWR VPWR
+ _02934_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_142_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 rvsingle.dp.rf.rf\[28\]\[9\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold611 rvsingle.dp.rf.rf\[13\]\[17\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold622 rvsingle.dp.rf.rf\[30\]\[7\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold633 rvsingle.dp.rf.rf\[16\]\[4\] VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold644 rvsingle.dp.rf.rf\[31\]\[9\] VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold655 rvsingle.dp.rf.rf\[4\]\[15\] VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold666 rvsingle.dp.rf.rf\[8\]\[21\] VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold677 rvsingle.dp.rf.rf\[8\]\[13\] VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 rvsingle.dp.rf.rf\[30\]\[15\] VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 rvsingle.dp.rf.rf\[7\]\[30\] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _04781_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__buf_2
X_08915_ _01138_ rvsingle.dp.rf.rf\[28\]\[25\] VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__nor2_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ Instr[11] VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__clkbuf_4
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _03766_ _02100_ _02015_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08777_ _03697_ _01537_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__nand2_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ rvsingle.dp.rf.rf\[23\]\[5\] _02627_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__and2b_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07659_ _01191_ rvsingle.dp.rf.rf\[6\]\[5\] _01299_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10670_ _04755_ net454 _05235_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09329_ _01169_ _02259_ _01170_ _01063_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__o31a_2
XFILLER_0_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12340_ _04845_ net716 _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12271_ _04839_ net316 _06073_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11222_ _05295_ rvsingle.dp.rf.rf\[29\]\[19\] _05541_ VGND VGND VPWR VPWR _05550_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11153_ _05512_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__clkbuf_1
X_10104_ _02908_ DataAdr[30] _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__a21oi_1
X_11084_ _05477_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__clkbuf_1
X_10035_ _04841_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ _05939_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__buf_6
XFILLER_0_129_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10937_ _04824_ net349 _05387_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_971 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10868_ _04858_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12607_ clknet_leaf_0_clk _00065_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10799_ _05309_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12538_ clknet_leaf_4_clk _01022_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12469_ clknet_leaf_27_clk _00953_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06961_ rvsingle.dp.rf.rf\[27\]\[22\] _01865_ _01881_ VGND VGND VPWR VPWR _01882_
+ sky130_fd_sc_hd__o21ai_1
X_08700_ _01137_ rvsingle.dp.rf.rf\[10\]\[14\] VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__nor2_1
X_09680_ _04520_ _04453_ _04525_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[13\] sky130_fd_sc_hd__o21ai_1
X_06892_ rvsingle.dp.rf.rf\[0\]\[23\] rvsingle.dp.rf.rf\[1\]\[23\] rvsingle.dp.rf.rf\[2\]\[23\]
+ rvsingle.dp.rf.rf\[3\]\[23\] _01469_ _01471_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08631_ rvsingle.dp.rf.rf\[31\]\[12\] _01677_ _03551_ VGND VGND VPWR VPWR _03552_
+ sky130_fd_sc_hd__o21ai_1
X_08562_ _01184_ _03455_ _03482_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07513_ _01349_ rvsingle.dp.rf.rf\[10\]\[6\] VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08493_ _01544_ rvsingle.dp.rf.rf\[28\]\[13\] _01610_ VGND VGND VPWR VPWR _03414_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07444_ _02117_ rvsingle.dp.rf.rf\[16\]\[7\] VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07375_ rvsingle.dp.rf.rf\[27\]\[7\] _01424_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09114_ _01126_ rvsingle.dp.rf.rf\[22\]\[26\] _01605_ VGND VGND VPWR VPWR _04034_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06326_ _01189_ _01220_ _01239_ _01248_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__o211a_2
XFILLER_0_127_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09045_ _03857_ rvsingle.dp.rf.rf\[7\]\[27\] _01106_ _03964_ VGND VGND VPWR VPWR
+ _03965_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06257_ _01179_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold430 rvsingle.dp.rf.rf\[21\]\[28\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
X_06188_ _01111_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__clkbuf_8
Xhold441 rvsingle.dp.rf.rf\[19\]\[27\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 rvsingle.dp.rf.rf\[10\]\[30\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 rvsingle.dp.rf.rf\[20\]\[22\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold474 rvsingle.dp.rf.rf\[5\]\[30\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 rvsingle.dp.rf.rf\[20\]\[17\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold496 rvsingle.dp.rf.rf\[25\]\[25\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09947_ DataAdr[6] ReadData[6] _04751_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _04618_ PC[31] VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__nor2_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _01153_ _03110_ _03087_ _01178_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__a31o_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _05881_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__clkbuf_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_146_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_146_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11771_ _05748_ _05847_ _05840_ net95 VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _04892_ net430 _05257_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__mux2_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10653_ _05227_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13372_ clknet_leaf_148_clk _00800_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10584_ _05188_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12323_ _04801_ net593 _06110_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12254_ _04781_ rvsingle.dp.rf.rf\[5\]\[9\] _06074_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11205_ _05527_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__buf_8
XFILLER_0_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12185_ _05757_ net307 _06048_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__mux2_1
X_11136_ _05503_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__clkbuf_1
X_11067_ _05468_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__clkbuf_1
X_10018_ _04826_ _04575_ _04743_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__mux2_4
XFILLER_0_92_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_137_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_137_clk sky130_fd_sc_hd__clkbuf_16
X_11969_ _05951_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07160_ _01223_ _02074_ _02080_ _01317_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07091_ _01960_ _01075_ _01961_ _02011_ _01587_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09801_ _04627_ _04552_ _04631_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07993_ _01067_ _01078_ _01080_ _01099_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__o211ai_2
X_09732_ _04571_ _04572_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__nand2_1
X_06944_ _01087_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__buf_4
X_09663_ PC[12] _04508_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__nor2_1
X_06875_ _01645_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__buf_4
X_08614_ _01620_ _03531_ _03532_ _01131_ _03534_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09594_ _04367_ _04443_ _04444_ _04446_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[6\]
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08545_ _01229_ _03460_ _03462_ _03465_ _02438_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__o221ai_4
Xclkbuf_leaf_128_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_128_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08476_ _03389_ _03396_ _02315_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__nand3_2
XFILLER_0_77_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07427_ _02297_ _01656_ _01620_ _02347_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07358_ _01420_ rvsingle.dp.rf.rf\[10\]\[7\] _01300_ _02278_ VGND VGND VPWR VPWR
+ _02279_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_116_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06309_ _01231_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__clkbuf_4
X_07289_ _01317_ _02205_ _02209_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__nand3_2
XFILLER_0_103_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09028_ _03945_ _03782_ _03947_ _01506_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold260 rvsingle.dp.rf.rf\[6\]\[25\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 rvsingle.dp.rf.rf\[18\]\[23\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 rvsingle.dp.rf.rf\[12\]\[17\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 rvsingle.dp.rf.rf\[4\]\[25\] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ clknet_leaf_42_clk _00399_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ clknet_leaf_106_clk _00330_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_100 _01097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _01335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _01452_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_133 _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11823_ _05872_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__clkbuf_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_119_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _01567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_166 _01695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _01763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _05840_ net37 _05734_ _05841_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__a22o_1
XANTENNA_199 _04383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _04840_ net548 _05246_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__mux2_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11685_ _05801_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10636_ _05218_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13355_ clknet_leaf_86_clk _00783_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10567_ _04859_ rvsingle.dp.rf.rf\[9\]\[23\] _05151_ VGND VGND VPWR VPWR _05179_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12306_ _04764_ net481 _06099_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__mux2_1
X_13286_ clknet_leaf_122_clk _00744_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10498_ _04892_ _05099_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__nand2_1
X_12237_ _04718_ _06070_ _06071_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__a21oi_1
X_12168_ _05744_ net224 _06049_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__mux2_1
X_11119_ _05377_ net633 _05490_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__mux2_1
X_12099_ _06009_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__buf_6
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06660_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06591_ _01511_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08330_ _01267_ rvsingle.dp.rf.rf\[4\]\[8\] VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08261_ _03176_ _02527_ _03181_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__nand3_1
XFILLER_0_144_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07212_ rvsingle.dp.rf.rf\[15\]\[17\] _01861_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08192_ rvsingle.dp.rf.rf\[4\]\[11\] rvsingle.dp.rf.rf\[5\]\[11\] rvsingle.dp.rf.rf\[6\]\[11\]
+ rvsingle.dp.rf.rf\[7\]\[11\] _01426_ _01433_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07143_ _02046_ _02051_ _01593_ _02063_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_160_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07074_ rvsingle.dp.rf.rf\[13\]\[19\] _01630_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__and2b_1
XFILLER_0_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07976_ rvsingle.dp.rf.rf\[17\]\[0\] _01677_ _02485_ VGND VGND VPWR VPWR _02897_
+ sky130_fd_sc_hd__o21ai_1
X_09715_ _04553_ _04453_ _04557_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[16\] sky130_fd_sc_hd__o21ai_1
X_06927_ _01847_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__clkbuf_8
X_09646_ PC[11] _04493_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__and2_1
X_06858_ _01095_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__buf_6
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _04397_ PC[3] PC[4] _04429_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ rvsingle.dp.rf.rf\[7\]\[20\] _01688_ _01709_ VGND VGND VPWR VPWR _01710_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08528_ _01753_ rvsingle.dp.rf.rf\[6\]\[13\] _01596_ _03448_ VGND VGND VPWR VPWR
+ _03449_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08459_ _03377_ _02291_ _03379_ _01446_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_163_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11470_ _05686_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10421_ _04892_ net236 _05082_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13140_ clknet_leaf_58_clk _00598_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10352_ _05053_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13071_ clknet_leaf_27_clk _00529_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10283_ _04904_ net272 _05001_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__mux2_1
X_12022_ _05979_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12924_ clknet_leaf_148_clk _00382_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12855_ clknet_leaf_6_clk _00313_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _05724_ net298 _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__mux2_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ clknet_leaf_56_clk _00244_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _05769_ _05770_ _05792_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11668_ _05790_ _05772_ _05791_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13407_ clknet_leaf_1_clk _00835_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10619_ _04800_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__buf_2
XFILLER_0_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11599_ net185 _05726_ _05760_ _05737_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13338_ clknet_leaf_77_clk rvsingle.dp.PCNext\[15\] _00015_ VGND VGND VPWR VPWR PC[15]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13269_ clknet_leaf_24_clk _00727_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07830_ _02469_ _02696_ _02747_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__o22ai_4
X_07761_ _02672_ _02674_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_155_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09500_ _04377_ _03194_ _03217_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__and3_4
X_06712_ _01629_ _01631_ _01632_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07692_ _01847_ rvsingle.dp.rf.rf\[8\]\[5\] _02612_ _01667_ VGND VGND VPWR VPWR _02613_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09431_ _03047_ _03052_ _02967_ _03049_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__o211a_1
X_06643_ _01130_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__buf_8
XFILLER_0_149_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09362_ _04275_ _04277_ _04213_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__o21bai_2
X_06574_ _01488_ rvsingle.dp.rf.rf\[27\]\[21\] _01491_ _01494_ VGND VGND VPWR VPWR
+ _01495_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08313_ rvsingle.dp.rf.rf\[15\]\[8\] _01508_ _02059_ VGND VGND VPWR VPWR _03234_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09293_ _04169_ _04168_ _04137_ _04172_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_75_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_11 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_22 Instr[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_33 Instr[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08244_ _01191_ rvsingle.dp.rf.rf\[0\]\[10\] VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_44 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_55 ReadData[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_66 ReadData[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_77 ReadData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08175_ rvsingle.dp.rf.rf\[3\]\[11\] _01566_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__or2b_1
XANTENNA_88 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 ReadData[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07126_ rvsingle.dp.rf.rf\[3\]\[18\] _01567_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__or2b_1
X_07057_ _01655_ _01974_ _01975_ _01768_ _01977_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_30_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07959_ rvsingle.dp.rf.rf\[15\]\[0\] _02478_ _01490_ VGND VGND VPWR VPWR _02880_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10970_ _05364_ _05365_ _05368_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09629_ _04474_ _04453_ _04478_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[9\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12640_ clknet_leaf_118_clk _00098_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12571_ clknet_leaf_136_clk _01055_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11522_ _05713_ net395 _05706_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11453_ _05359_ net465 _05668_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10404_ _05063_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11384_ _05266_ net459 _05629_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13123_ clknet_leaf_123_clk _00581_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10335_ _04846_ net366 _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ clknet_leaf_134_clk _00512_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10266_ _05004_ _05007_ _04978_ net154 VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__a2bb2o_1
X_12005_ _05716_ net239 _05960_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__mux2_1
X_10197_ _04904_ net301 _04952_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12907_ clknet_leaf_88_clk _00365_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12838_ clknet_leaf_113_clk _00296_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12769_ clknet_leaf_141_clk _00227_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06290_ rvsingle.dp.rf.rf\[0\]\[30\] rvsingle.dp.rf.rf\[1\]\[30\] rvsingle.dp.rf.rf\[2\]\[30\]
+ rvsingle.dp.rf.rf\[3\]\[30\] _01196_ _01203_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold804 rvsingle.dp.rf.rf\[30\]\[14\] VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold815 rvsingle.dp.rf.rf\[31\]\[11\] VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09980_ _04794_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08931_ rvsingle.dp.rf.rf\[17\]\[25\] _03839_ _01497_ _03851_ VGND VGND VPWR VPWR
+ _03852_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08862_ _03777_ _03780_ _03781_ _03782_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__o2bb2ai_1
X_07813_ _01797_ rvsingle.dp.rf.rf\[22\]\[3\] VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__nor2_1
X_08793_ rvsingle.dp.rf.rf\[12\]\[15\] rvsingle.dp.rf.rf\[13\]\[15\] rvsingle.dp.rf.rf\[14\]\[15\]
+ rvsingle.dp.rf.rf\[15\]\[15\] _01335_ _01199_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__mux4_2
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07744_ _02315_ _02593_ _02607_ _01246_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07675_ _01327_ rvsingle.dp.rf.rf\[30\]\[5\] VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09414_ _03064_ _04295_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__nand2_1
X_06626_ rvsingle.dp.rf.rf\[13\]\[21\] _01540_ _01543_ _01546_ VGND VGND VPWR VPWR
+ _01547_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_59_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09345_ net820 _03483_ _03572_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06557_ _01446_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09276_ _03909_ _03827_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06488_ _01408_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08227_ rvsingle.dp.rf.rf\[28\]\[10\] rvsingle.dp.rf.rf\[29\]\[10\] rvsingle.dp.rf.rf\[30\]\[10\]
+ rvsingle.dp.rf.rf\[31\]\[10\] _02450_ _01708_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08158_ rvsingle.dp.rf.rf\[27\]\[11\] _01566_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__or2b_1
XFILLER_0_133_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07109_ _01566_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__buf_8
X_08089_ _01642_ rvsingle.dp.rf.rf\[8\]\[1\] VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10120_ _04722_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__buf_4
XFILLER_0_101_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_99_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
X_10051_ _04140_ _04141_ _04732_ ReadData[23] VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__or4b_1
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10953_ _05404_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10884_ _05361_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12623_ clknet_leaf_36_clk _00081_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12554_ clknet_leaf_84_clk _01038_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11505_ _05704_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12485_ clknet_leaf_114_clk _00969_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11436_ _05398_ net801 _05657_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11367_ _05606_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__buf_8
XFILLER_0_132_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13106_ clknet_leaf_56_clk _00564_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _04802_ net733 _05033_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _05400_ rvsingle.dp.rf.rf\[15\]\[21\] _05591_ VGND VGND VPWR VPWR _05592_
+ sky130_fd_sc_hd__mux2_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ clknet_leaf_44_clk _00495_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _04997_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07460_ _02030_ rvsingle.dp.rf.rf\[24\]\[6\] VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06411_ _01326_ _01311_ _01209_ _01332_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07391_ rvsingle.dp.rf.rf\[23\]\[7\] _01827_ _02311_ VGND VGND VPWR VPWR _02312_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
X_09130_ _01153_ _04031_ _04049_ _01482_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__nand4_1
X_06342_ _01138_ rvsingle.dp.rf.rf\[12\]\[29\] VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09061_ _01180_ _03980_ _01184_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__o21a_2
XFILLER_0_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06273_ _01195_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08012_ _01327_ rvsingle.dp.rf.rf\[20\]\[0\] VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold601 rvsingle.dp.rf.rf\[26\]\[12\] VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold612 rvsingle.dp.rf.rf\[28\]\[12\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold623 rvsingle.dp.rf.rf\[12\]\[4\] VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 rvsingle.dp.rf.rf\[18\]\[21\] VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold645 rvsingle.dp.rf.rf\[13\]\[26\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 rvsingle.dp.rf.rf\[28\]\[6\] VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 rvsingle.dp.rf.rf\[3\]\[29\] VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 rvsingle.dp.rf.rf\[24\]\[25\] VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ _04780_ _04477_ _04743_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__mux2_4
Xhold689 rvsingle.dp.rf.rf\[31\]\[2\] VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ _01257_ rvsingle.dp.rf.rf\[24\]\[25\] _03834_ _01856_ VGND VGND VPWR VPWR
+ _03835_ sky130_fd_sc_hd__o211a_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__clkbuf_2
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _02012_ _02014_ _01959_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__a21oi_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08776_ _01962_ _01128_ _03673_ _03696_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__o211ai_4
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ _01769_ rvsingle.dp.rf.rf\[22\]\[5\] _01104_ VGND VGND VPWR VPWR _02648_
+ sky130_fd_sc_hd__o21ai_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07658_ rvsingle.dp.rf.rf\[5\]\[5\] _02271_ _02268_ _02578_ VGND VGND VPWR VPWR _02579_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06609_ _01103_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
X_07589_ _02506_ _02507_ _02509_ _01600_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_137_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09328_ _01581_ _03879_ _01066_ _01075_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09259_ _03983_ _04053_ _04056_ _04057_ _03982_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12270_ _06085_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11221_ _05549_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11152_ _05295_ net673 _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__mux2_1
X_10103_ _04879_ _04880_ _04881_ ReadData[30] _04715_ VGND VGND VPWR VPWR _04900_
+ sky130_fd_sc_hd__o311a_1
X_11083_ _05476_ net290 _05469_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__mux2_1
X_10034_ _04840_ net437 _04791_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__mux2_1
X_11985_ _05959_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10936_ _05394_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10867_ _04853_ _05183_ _05336_ _05351_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ clknet_leaf_150_clk _00064_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10798_ _04892_ net344 _05298_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__mux2_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12537_ clknet_leaf_7_clk _01021_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12468_ clknet_leaf_20_clk _00952_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11419_ _05658_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12399_ clknet_leaf_36_clk _00883_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06960_ _01558_ rvsingle.dp.rf.rf\[26\]\[22\] _01880_ VGND VGND VPWR VPWR _01881_
+ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_3_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_06891_ _01208_ _01805_ _01811_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08630_ _01561_ rvsingle.dp.rf.rf\[30\]\[12\] _01530_ VGND VGND VPWR VPWR _03551_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08561_ _01201_ _01351_ _03467_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_49_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07512_ rvsingle.dp.rf.rf\[8\]\[6\] rvsingle.dp.rf.rf\[9\]\[6\] _01730_ VGND VGND
+ VPWR VPWR _02433_ sky130_fd_sc_hd__mux2_1
X_08492_ rvsingle.dp.rf.rf\[31\]\[13\] _01087_ _01880_ VGND VGND VPWR VPWR _03413_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07443_ _01155_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__buf_6
XFILLER_0_71_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07374_ _01192_ rvsingle.dp.rf.rf\[26\]\[7\] _01199_ VGND VGND VPWR VPWR _02295_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09113_ _03839_ rvsingle.dp.rf.rf\[21\]\[26\] _04032_ VGND VGND VPWR VPWR _04033_
+ sky130_fd_sc_hd__o21ai_1
X_06325_ _01247_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09044_ _01744_ rvsingle.dp.rf.rf\[6\]\[27\] VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__or2_1
X_06256_ _01171_ _01176_ _01178_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold420 rvsingle.dp.rf.rf\[2\]\[24\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 rvsingle.dp.rf.rf\[29\]\[10\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ _01110_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__buf_8
Xhold442 rvsingle.dp.rf.rf\[11\]\[28\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 rvsingle.dp.rf.rf\[24\]\[27\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 rvsingle.dp.rf.rf\[28\]\[22\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 rvsingle.dp.rf.rf\[30\]\[25\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 rvsingle.dp.rf.rf\[11\]\[23\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 rvsingle.dp.rf.rf\[7\]\[27\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
X_09946_ _01169_ _02259_ _01170_ _04445_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__or4b_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _04693_ _04694_ _04696_ _04697_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__a22oi_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _03313_ _03405_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__a21oi_1
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ rvsingle.dp.rf.rf\[15\]\[15\] _01508_ _02059_ VGND VGND VPWR VPWR _03680_
+ sky130_fd_sc_hd__o21ai_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _05747_ _05847_ _05840_ net165 VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _05264_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10652_ _04892_ net330 _05219_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13371_ clknet_leaf_138_clk _00799_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10583_ _05187_ net334 _05151_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12322_ _06112_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12253_ _06079_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__clkbuf_1
X_11204_ _05540_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12184_ _04853_ _05766_ _05336_ _06058_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__a31o_1
X_11135_ _05334_ net432 _05499_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11066_ _05428_ net448 _05460_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__mux2_1
X_10017_ DataAdr[18] ReadData[18] _04750_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11968_ _04785_ net560 _05949_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10919_ _05384_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__clkbuf_1
X_11899_ _05901_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__buf_6
XFILLER_0_156_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07090_ _01962_ _01128_ _01985_ _02010_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09800_ _04628_ _04631_ _04634_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__a21o_1
X_07992_ _01175_ net823 Instr[7] _02912_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06943_ _01861_ rvsingle.dp.rf.rf\[7\]\[22\] _01655_ _01863_ VGND VGND VPWR VPWR
+ _01864_ sky130_fd_sc_hd__o211ai_1
X_09731_ _01224_ _02912_ _04506_ _04507_ PC[18] VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__a311o_1
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09662_ _04508_ PC[12] VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__and2_1
X_06874_ rvsingle.dp.rf.rf\[23\]\[23\] _01097_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__and2b_1
X_08613_ _01382_ rvsingle.dp.rf.rf\[2\]\[12\] _01777_ _03533_ VGND VGND VPWR VPWR
+ _03534_ sky130_fd_sc_hd__o211ai_1
X_09593_ _04422_ _04423_ _04445_ _04427_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _03464_ _02291_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08475_ _01207_ _03390_ _03395_ _02447_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07426_ _01567_ rvsingle.dp.rf.rf\[24\]\[7\] VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07357_ rvsingle.dp.rf.rf\[11\]\[7\] _02163_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06308_ _01230_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07288_ _02191_ _02206_ _02208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09027_ rvsingle.dp.rf.rf\[23\]\[27\] _01089_ _03946_ VGND VGND VPWR VPWR _03947_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06239_ _01090_ rvsingle.dp.rf.rf\[31\]\[30\] _01107_ _01162_ VGND VGND VPWR VPWR
+ _01163_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold250 rvsingle.dp.rf.rf\[19\]\[23\] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold261 rvsingle.dp.rf.rf\[30\]\[29\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold272 rvsingle.dp.rf.rf\[27\]\[30\] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 rvsingle.dp.rf.rf\[26\]\[9\] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 rvsingle.dp.rf.rf\[9\]\[28\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
X_09929_ _04425_ _04752_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12940_ clknet_leaf_52_clk _00398_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ clknet_leaf_99_clk _00329_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _01148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _01420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _01487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_134 _01520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11822_ _05428_ net269 _05863_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__mux2_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _01567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _01695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_178 _01769_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11753_ _05830_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__buf_6
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_189 _02011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10704_ _05255_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11684_ _05496_ net719 _05795_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10635_ _04840_ net609 _05205_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13354_ clknet_leaf_80_clk rvsingle.dp.PCNext\[31\] _00031_ VGND VGND VPWR VPWR PC[31]
+ sky130_fd_sc_hd__dfrtp_4
X_10566_ net27 _05155_ _05178_ _05157_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12305_ _06103_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13285_ clknet_leaf_124_clk _00743_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10497_ _05136_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12236_ _05145_ _05830_ net164 VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12167_ net85 _06049_ _06021_ _04985_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__a22o_1
X_11118_ _05493_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__clkbuf_1
X_12098_ _06018_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__clkbuf_1
X_11049_ _04919_ _04733_ _05371_ _04737_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__or4b_2
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06590_ _01110_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__buf_8
XFILLER_0_87_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08260_ _01092_ _03177_ _03178_ _01511_ _03180_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_157_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07211_ _01744_ rvsingle.dp.rf.rf\[14\]\[17\] _01648_ VGND VGND VPWR VPWR _02132_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08191_ _02473_ _02318_ _01961_ _03111_ _01580_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07142_ _02056_ _02062_ _01506_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__nand3_1
XFILLER_0_171_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07073_ _01518_ rvsingle.dp.rf.rf\[12\]\[19\] _01611_ VGND VGND VPWR VPWR _01994_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07975_ rvsingle.dp.rf.rf\[16\]\[0\] _01603_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__nor2_1
X_09714_ _04454_ _04455_ _04556_ _04459_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__o211ai_1
X_06926_ _01752_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__buf_6
X_06857_ _01656_ rvsingle.dp.rf.rf\[24\]\[23\] _01777_ VGND VGND VPWR VPWR _01778_
+ sky130_fd_sc_hd__o21bai_1
X_09645_ _04492_ Instr[31] _04369_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__mux2_2
XFILLER_0_93_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09576_ _04429_ _04421_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _01707_ rvsingle.dp.rf.rf\[6\]\[20\] _01708_ VGND VGND VPWR VPWR _01709_
+ sky130_fd_sc_hd__o21a_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ rvsingle.dp.rf.rf\[7\]\[13\] _01752_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08458_ rvsingle.dp.rf.rf\[7\]\[9\] _01295_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07409_ rvsingle.dp.rf.rf\[11\]\[7\] _01557_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08389_ _03301_ _03303_ _03309_ _02315_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10420_ _05091_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10351_ _04898_ net446 _05044_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13070_ clknet_leaf_52_clk _00528_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10282_ _05015_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
X_12021_ _05531_ rvsingle.dp.rf.rf\[8\]\[3\] _05976_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__mux2_1
X_12923_ clknet_leaf_141_clk _00381_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12854_ clknet_leaf_34_clk _00312_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _05862_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__buf_6
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ clknet_leaf_56_clk _00243_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11736_ net48 VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11667_ _05769_ _05770_ _05772_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13406_ clknet_leaf_0_clk _00834_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10618_ _05208_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__clkbuf_1
X_11598_ _04869_ _04968_ _04967_ _05097_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10549_ _05167_ _05169_ _05155_ net139 VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__a2bb2o_1
X_13337_ clknet_leaf_75_clk rvsingle.dp.PCNext\[14\] _00014_ VGND VGND VPWR VPWR PC[14]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13268_ clknet_leaf_58_clk _00726_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12219_ _06068_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__inv_2
X_13199_ clknet_leaf_44_clk _00657_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07760_ _01711_ _02675_ _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__o21ai_1
X_06711_ _01110_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07691_ rvsingle.dp.rf.rf\[9\]\[5\] _01752_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__or2b_1
XFILLER_0_91_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09430_ _03047_ _03052_ _03049_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__o21ai_1
X_06642_ rvsingle.dp.rf.rf\[1\]\[21\] _01562_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09361_ _03765_ _04276_ _04214_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__a21oi_2
X_06573_ _01493_ rvsingle.dp.rf.rf\[26\]\[21\] VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08312_ _01513_ rvsingle.dp.rf.rf\[14\]\[8\] VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09292_ _01925_ _01928_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 Instr[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08243_ rvsingle.dp.rf.rf\[3\]\[10\] _01827_ _01808_ VGND VGND VPWR VPWR _03164_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_34 Instr[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_45 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_56 ReadData[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 ReadData[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_78 ReadData[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08174_ _03093_ _03094_ _01110_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_160_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_89 ReadData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07125_ _02042_ _02043_ _02045_ _01112_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07056_ _01256_ rvsingle.dp.rf.rf\[26\]\[19\] _01660_ _01976_ VGND VGND VPWR VPWR
+ _01977_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_88_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07958_ rvsingle.dp.rf.rf\[14\]\[0\] _01518_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06909_ _01827_ rvsingle.dp.rf.rf\[27\]\[23\] _01808_ _01829_ VGND VGND VPWR VPWR
+ _01830_ sky130_fd_sc_hd__o211a_1
X_07889_ rvsingle.dp.rf.rf\[9\]\[2\] _02288_ _01308_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09628_ _04454_ _04455_ _04477_ _04459_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_97_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09559_ Instr[11] _01078_ PC[4] _02531_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12570_ clknet_leaf_5_clk _01054_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11521_ _04885_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__buf_2
XFILLER_0_53_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11452_ _05675_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10403_ _05083_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__clkbuf_1
X_11383_ _05637_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13122_ clknet_leaf_136_clk _00580_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10334_ _05021_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__buf_6
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ clknet_leaf_143_clk _00511_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10265_ _04846_ _04970_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__nand2_1
X_12004_ _05137_ _05847_ _05940_ net252 VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__a2bb2o_1
X_10196_ _04961_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12906_ clknet_leaf_95_clk _00364_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12837_ clknet_leaf_113_clk _00295_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ clknet_leaf_117_clk _00226_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11719_ _05819_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__clkbuf_1
X_12699_ clknet_leaf_137_clk _00157_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold805 rvsingle.dp.rf.rf\[29\]\[2\] VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold816 rvsingle.dp.rf.rf\[29\]\[3\] VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08930_ _01562_ rvsingle.dp.rf.rf\[16\]\[25\] VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08861_ _01632_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__buf_4
X_07812_ rvsingle.dp.rf.rf\[23\]\[3\] VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__inv_2
X_08792_ _03705_ _03712_ _02315_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__nand3_4
X_07743_ Instr[25] _01537_ _01183_ _02663_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__o211ai_2
X_07674_ rvsingle.dp.rf.rf\[28\]\[5\] rvsingle.dp.rf.rf\[29\]\[5\] _01419_ VGND VGND
+ VPWR VPWR _02595_ sky130_fd_sc_hd__mux2_1
X_06625_ _01545_ rvsingle.dp.rf.rf\[12\]\[21\] VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__or2_1
X_09413_ _02263_ _04323_ _04324_ VGND VGND VPWR VPWR DataAdr[16] sky130_fd_sc_hd__o21ai_4
XFILLER_0_88_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06556_ _01476_ _01445_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__nand2_1
X_09344_ _04258_ _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__nor2_2
XFILLER_0_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09275_ _04051_ _04052_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06487_ _01375_ _01406_ _01407_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08226_ _02302_ _03146_ _02447_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08157_ _03076_ _03077_ _01564_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07108_ rvsingle.dp.rf.rf\[17\]\[18\] _01088_ _01668_ VGND VGND VPWR VPWR _02029_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08088_ rvsingle.dp.rf.rf\[11\]\[1\] _01645_ _01647_ VGND VGND VPWR VPWR _03009_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07039_ _01064_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__buf_8
XFILLER_0_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10050_ _04854_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10952_ _05352_ net271 _05401_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10883_ _05266_ rvsingle.dp.rf.rf\[1\]\[29\] _05319_ VGND VGND VPWR VPWR _05361_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12622_ clknet_leaf_71_clk _00080_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12553_ clknet_leaf_96_clk _01037_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11504_ _05295_ net695 _05695_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12484_ clknet_leaf_109_clk _00968_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11435_ _05666_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11366_ _05628_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__clkbuf_1
X_10317_ _05035_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__clkbuf_1
X_13105_ clknet_leaf_57_clk _00563_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _05568_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__buf_6
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13036_ clknet_leaf_50_clk _00494_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _04808_ rvsingle.dp.rf.rf\[27\]\[14\] _04989_ VGND VGND VPWR VPWR _04997_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10179_ _04846_ net279 _04952_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06410_ _01297_ rvsingle.dp.rf.rf\[31\]\[29\] _01201_ _01331_ VGND VGND VPWR VPWR
+ _01332_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07390_ _01725_ rvsingle.dp.rf.rf\[22\]\[7\] _01198_ VGND VGND VPWR VPWR _02311_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06341_ rvsingle.dp.rf.rf\[8\]\[29\] rvsingle.dp.rf.rf\[9\]\[29\] rvsingle.dp.rf.rf\[10\]\[29\]
+ rvsingle.dp.rf.rf\[11\]\[29\] _01127_ _01261_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09060_ _01153_ _03956_ _03977_ _01084_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__and4_1
X_06272_ _01194_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08011_ _02927_ _02928_ _01206_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold602 rvsingle.dp.rf.rf\[2\]\[14\] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold613 rvsingle.dp.rf.rf\[8\]\[10\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 rvsingle.dp.rf.rf\[22\]\[29\] VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold635 rvsingle.dp.rf.rf\[23\]\[22\] VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold646 rvsingle.dp.rf.rf\[15\]\[6\] VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 rvsingle.dp.rf.rf\[31\]\[27\] VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold668 rvsingle.dp.rf.rf\[29\]\[17\] VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 rvsingle.dp.rf.rf\[4\]\[5\] VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ DataAdr[9] ReadData[9] _04750_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08913_ rvsingle.dp.rf.rf\[25\]\[25\] _01126_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__or2b_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _04713_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__buf_2
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _02181_ _03762_ _03764_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__o21ai_4
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _01593_ _03684_ _03695_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__nand3_4
XFILLER_0_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _02645_ _01780_ _02337_ _02646_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__a211oi_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07657_ _01690_ rvsingle.dp.rf.rf\[4\]\[5\] VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__or2_1
X_06608_ rvsingle.dp.rf.rf\[17\]\[21\] _01509_ _01497_ VGND VGND VPWR VPWR _01529_
+ sky130_fd_sc_hd__o21ai_1
X_07588_ _01513_ rvsingle.dp.rf.rf\[16\]\[4\] _02508_ _01496_ VGND VGND VPWR VPWR
+ _02509_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_168_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09327_ _03830_ _04238_ _04240_ _03827_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06539_ _01206_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09258_ _03775_ _03910_ _04056_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__nand3_1
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08209_ rvsingle.dp.rf.rf\[16\]\[11\] rvsingle.dp.rf.rf\[17\]\[11\] rvsingle.dp.rf.rf\[18\]\[11\]
+ rvsingle.dp.rf.rf\[19\]\[11\] _01416_ _01300_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09189_ _04102_ _01118_ _01147_ _04108_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__a211o_1
XFILLER_0_160_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11220_ _05439_ rvsingle.dp.rf.rf\[29\]\[18\] _05541_ VGND VGND VPWR VPWR _05549_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11151_ _05489_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__buf_8
XFILLER_0_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10102_ _04899_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
X_11082_ _04823_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__buf_2
XFILLER_0_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10033_ _04839_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__clkbuf_4
X_11984_ _05173_ net327 _05949_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10935_ _05291_ rvsingle.dp.rf.rf\[18\]\[16\] _05387_ VGND VGND VPWR VPWR _05394_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10866_ _05337_ _05338_ _05339_ _05084_ net206 VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__o41a_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12605_ clknet_leaf_143_clk _00063_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_995 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10797_ _05308_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12536_ clknet_leaf_34_clk _01020_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12467_ clknet_leaf_29_clk _00951_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11418_ _05334_ net640 _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__mux2_1
X_12398_ clknet_leaf_53_clk _00882_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11349_ _05207_ net776 _05618_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13019_ clknet_leaf_136_clk _00477_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_06890_ _01461_ _01807_ _01810_ _01218_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__a31oi_1
X_08560_ _01316_ _03473_ _03480_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__nand3_2
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07511_ _01065_ _02318_ _01178_ _02427_ _02431_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08491_ _01862_ rvsingle.dp.rf.rf\[30\]\[13\] VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07442_ _02361_ _02362_ _02323_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07373_ rvsingle.dp.rf.rf\[28\]\[7\] rvsingle.dp.rf.rf\[29\]\[7\] rvsingle.dp.rf.rf\[30\]\[7\]
+ rvsingle.dp.rf.rf\[31\]\[7\] _01426_ _01433_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__mux4_2
XFILLER_0_18_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09112_ _01126_ rvsingle.dp.rf.rf\[20\]\[26\] _01531_ VGND VGND VPWR VPWR _04032_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06324_ _01246_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__buf_8
XFILLER_0_33_807 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_894 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09043_ rvsingle.dp.rf.rf\[5\]\[27\] _03778_ _01093_ _03962_ VGND VGND VPWR VPWR
+ _03963_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06255_ net822 VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold410 rvsingle.dp.rf.rf\[14\]\[6\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
X_06186_ Instr[22] VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__clkbuf_8
Xhold421 rvsingle.dp.rf.rf\[28\]\[26\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 rvsingle.dp.rf.rf\[16\]\[11\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold443 rvsingle.dp.rf.rf\[31\]\[29\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 rvsingle.dp.rf.rf\[21\]\[3\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 rvsingle.dp.rf.rf\[13\]\[28\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 rvsingle.dp.rf.rf\[8\]\[18\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 rvsingle.dp.rf.rf\[6\]\[7\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 rvsingle.dp.rf.rf\[23\]\[13\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ _04766_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__clkbuf_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _04701_ _04698_ _04702_ _04703_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__nand4b_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _02469_ _03747_ _03404_ _03402_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__a2bb2oi_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _01513_ rvsingle.dp.rf.rf\[14\]\[15\] VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__nor2_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _01607_ rvsingle.dp.rf.rf\[2\]\[5\] _01596_ _02629_ VGND VGND VPWR VPWR _02630_
+ sky130_fd_sc_hd__o211ai_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ rvsingle.dp.rf.rf\[17\]\[14\] _01255_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__and2b_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10720_ _04886_ net750 _05257_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__mux2_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10651_ _05226_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13370_ clknet_leaf_14_clk _00798_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10582_ _04903_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__buf_2
XFILLER_0_51_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12321_ _04795_ net506 _06110_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12252_ _04777_ rvsingle.dp.rf.rf\[5\]\[8\] _06074_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11203_ _05385_ net431 _05528_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12183_ _05337_ _05338_ _05339_ _05003_ net207 VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__o41a_1
X_11134_ _05502_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__clkbuf_1
X_11065_ _05467_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__clkbuf_1
X_10016_ _04825_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11967_ _05950_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10918_ _04782_ net577 _05373_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11898_ _05912_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10849_ _04916_ _04918_ _04965_ _04807_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__or4b_2
XFILLER_0_6_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12519_ clknet_leaf_100_clk _01003_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07991_ _01076_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ _04570_ PC[18] VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__nand2_1
X_06942_ _01862_ rvsingle.dp.rf.rf\[6\]\[22\] VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09661_ Instr[12] _04505_ _04506_ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__a31o_1
X_06873_ _01562_ rvsingle.dp.rf.rf\[22\]\[23\] VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08612_ rvsingle.dp.rf.rf\[3\]\[12\] _01779_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__or2b_1
X_09592_ _04397_ PC[3] PC[4] _04429_ PC[6] VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__a41o_1
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08543_ rvsingle.dp.rf.rf\[29\]\[13\] _02275_ _01436_ _03463_ VGND VGND VPWR VPWR
+ _03464_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08474_ _03391_ _03392_ _02543_ _03394_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07425_ _01377_ _02333_ _02345_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__nand3_4
XFILLER_0_58_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07356_ _02275_ rvsingle.dp.rf.rf\[9\]\[7\] _02276_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06307_ _01229_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07287_ _01445_ _02207_ _01447_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__o21a_1
XFILLER_0_171_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09026_ _01098_ rvsingle.dp.rf.rf\[22\]\[27\] _01655_ VGND VGND VPWR VPWR _03946_
+ sky130_fd_sc_hd__o21a_1
X_06238_ _01139_ rvsingle.dp.rf.rf\[30\]\[30\] VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold240 rvsingle.dp.rf.rf\[6\]\[27\] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
X_06169_ _01092_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__buf_4
Xhold251 rvsingle.dp.rf.rf\[7\]\[12\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 rvsingle.dp.rf.rf\[4\]\[26\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 rvsingle.dp.rf.rf\[28\]\[20\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 rvsingle.dp.rf.rf\[30\]\[11\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 rvsingle.dp.rf.rf\[14\]\[30\] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ DataAdr[3] ReadData[3] _04751_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__mux2_1
X_09859_ _04686_ _04687_ _04685_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__a21o_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ clknet_leaf_108_clk _00328_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _01422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11821_ _05871_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__clkbuf_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _01492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 _01520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _01595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _01660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _01695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _05837_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__buf_4
XFILLER_0_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_179 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _04834_ rvsingle.dp.rf.rf\[21\]\[19\] _05246_ VGND VGND VPWR VPWR _05255_
+ sky130_fd_sc_hd__mux2_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11683_ _05800_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10634_ _05217_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13353_ clknet_leaf_80_clk rvsingle.dp.PCNext\[30\] _00030_ VGND VGND VPWR VPWR PC[30]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10565_ _04879_ _04881_ _04880_ _05058_ _04852_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__o311a_2
XFILLER_0_162_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12304_ _04759_ net706 _06099_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13284_ clknet_leaf_131_clk _00742_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10496_ _04886_ net453 _05126_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12235_ _04721_ _05058_ _05830_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__and3_1
X_12166_ net21 _06052_ _05332_ _04985_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__a22o_1
X_11117_ _04755_ net702 _05490_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__mux2_1
X_12097_ _05740_ net356 _06010_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__mux2_1
X_11048_ _05314_ _05456_ _05458_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12999_ clknet_leaf_98_clk _00457_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07210_ _01759_ _02129_ _02130_ _01768_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_7_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08190_ _01150_ _01139_ _03087_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07141_ _02057_ _02058_ _01565_ _02061_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_171_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07072_ _01991_ _01383_ _01992_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07974_ _01600_ _02892_ _02894_ _02364_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__a31o_1
X_09713_ _04554_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__nor2_2
X_06925_ _01841_ _01843_ _01844_ _01845_ _01112_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__o221a_1
X_09644_ Instr[7] _04140_ MemWrite _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__o31a_1
X_06856_ _01258_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__buf_8
XFILLER_0_69_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09575_ PC[5] VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__buf_2
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ _01454_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__buf_6
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ rvsingle.dp.rf.rf\[5\]\[13\] _01498_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__and2b_1
X_08457_ _01468_ rvsingle.dp.rf.rf\[6\]\[9\] _01198_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07408_ _01130_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__buf_4
XFILLER_0_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08388_ _01694_ _03304_ _03308_ _01699_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07339_ _02259_ _01173_ _01174_ _01169_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__nor4_2
XFILLER_0_122_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10350_ _05052_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09009_ rvsingle.dp.rf.rf\[12\]\[27\] rvsingle.dp.rf.rf\[13\]\[27\] rvsingle.dp.rf.rf\[14\]\[27\]
+ rvsingle.dp.rf.rf\[15\]\[27\] _01336_ _01200_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10281_ _04898_ net710 _05001_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _05978_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__clkbuf_1
X_12922_ clknet_leaf_3_clk _00380_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ clknet_leaf_37_clk _00311_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _04723_ _04928_ _04975_ _04722_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__or4b_4
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ clknet_leaf_68_clk _00242_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11735_ _05827_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__clkbuf_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ net51 VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13405_ clknet_leaf_143_clk _00833_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10617_ _05207_ rvsingle.dp.rf.rf\[22\]\[12\] _05205_ VGND VGND VPWR VPWR _05208_
+ sky130_fd_sc_hd__mux2_1
X_11597_ _05149_ _05759_ _05731_ net102 VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13336_ clknet_leaf_75_clk rvsingle.dp.PCNext\[13\] _00013_ VGND VGND VPWR VPWR PC[13]
+ sky130_fd_sc_hd__dfrtp_4
X_10548_ _04808_ _05144_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13267_ clknet_leaf_67_clk _00725_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10479_ _04834_ net625 _05126_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12218_ _06068_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13198_ clknet_leaf_53_clk _00656_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12149_ _05316_ _04973_ net28 VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__a21oi_1
X_06710_ rvsingle.dp.rf.rf\[7\]\[20\] _01630_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07690_ rvsingle.dp.rf.rf\[11\]\[5\] _01087_ _01654_ VGND VGND VPWR VPWR _02611_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06641_ _01561_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09360_ _04165_ _02184_ _02265_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__nand3_1
X_06572_ _01492_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__buf_8
XFILLER_0_164_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08311_ Instr[28] VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09291_ _04199_ _04201_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 DataAdr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08242_ _01726_ rvsingle.dp.rf.rf\[2\]\[10\] VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_24 Instr[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 Instr[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_46 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_57 ReadData[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_68 ReadData[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08173_ rvsingle.dp.rf.rf\[1\]\[11\] _01594_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_79 ReadData[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07124_ rvsingle.dp.rf.rf\[5\]\[18\] _01540_ _01759_ _02044_ VGND VGND VPWR VPWR
+ _02045_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_144_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07055_ rvsingle.dp.rf.rf\[27\]\[19\] _01650_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__or2b_1
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07957_ _02876_ _01643_ _01105_ _02877_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__a211oi_2
X_06908_ _01828_ rvsingle.dp.rf.rf\[26\]\[23\] VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07888_ _01726_ rvsingle.dp.rf.rf\[8\]\[2\] VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__nor2_1
X_09627_ _04475_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__nor2_1
X_06839_ _01603_ rvsingle.dp.rf.rf\[6\]\[23\] VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09558_ _04367_ _04406_ _04413_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[3\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08509_ _01382_ rvsingle.dp.rf.rf\[10\]\[13\] VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09489_ _04385_ VGND VGND VPWR VPWR WriteData[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11520_ _05712_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11451_ _05307_ rvsingle.dp.rf.rf\[13\]\[27\] _05668_ VGND VGND VPWR VPWR _05675_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10402_ _04828_ rvsingle.dp.rf.rf\[25\]\[18\] _05082_ VGND VGND VPWR VPWR _05083_
+ sky130_fd_sc_hd__mux2_1
X_11382_ _05359_ net427 _05629_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13121_ clknet_leaf_126_clk _00579_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10333_ _05043_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13052_ clknet_leaf_13_clk _00510_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10264_ net26 _04978_ _05006_ _04985_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12003_ _05968_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__clkbuf_1
X_10195_ _04898_ net306 _04952_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12905_ clknet_leaf_97_clk _00363_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12836_ clknet_leaf_101_clk _00294_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ clknet_leaf_3_clk _00225_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _05300_ net587 _05817_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12698_ clknet_leaf_15_clk _00156_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11649_ _05400_ net813 _05775_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold806 rvsingle.dp.rf.rf\[15\]\[8\] VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold817 rvsingle.dp.rf.rf\[18\]\[13\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ clknet_leaf_121_clk _00777_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08860_ rvsingle.dp.rf.rf\[16\]\[24\] rvsingle.dp.rf.rf\[17\]\[24\] rvsingle.dp.rf.rf\[18\]\[24\]
+ rvsingle.dp.rf.rf\[19\]\[24\] _01493_ _01612_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__mux4_1
X_07811_ _02726_ _02731_ _02491_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__nand3_1
X_08791_ _01461_ _03706_ _03711_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07742_ _02662_ _01481_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07673_ rvsingle.dp.rf.rf\[24\]\[5\] rvsingle.dp.rf.rf\[25\]\[5\] rvsingle.dp.rf.rf\[26\]\[5\]
+ rvsingle.dp.rf.rf\[27\]\[5\] _01328_ _01455_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__mux4_1
X_09412_ _02265_ _04165_ _04247_ _04117_ _04251_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__o2111ai_4
X_06624_ _01544_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09343_ _03064_ _04148_ _04161_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__a21oi_1
X_06555_ rvsingle.dp.rf.rf\[13\]\[21\] _01441_ _01437_ _01475_ VGND VGND VPWR VPWR
+ _01476_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_90_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09274_ DataAdr[29] DataAdr[30] VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__nor2_1
X_06486_ _01085_ WriteData[28] _01180_ _01184_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08225_ rvsingle.dp.rf.rf\[16\]\[10\] rvsingle.dp.rf.rf\[17\]\[10\] rvsingle.dp.rf.rf\[18\]\[10\]
+ rvsingle.dp.rf.rf\[19\]\[10\] _01328_ _01455_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08156_ rvsingle.dp.rf.rf\[25\]\[11\] _01492_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07107_ _01666_ rvsingle.dp.rf.rf\[16\]\[18\] VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08087_ _01797_ rvsingle.dp.rf.rf\[10\]\[1\] VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07038_ _01247_ _01942_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08989_ _03907_ _03880_ _03881_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__or3_2
XFILLER_0_98_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10951_ _05403_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10882_ _05360_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12621_ clknet_leaf_43_clk _00079_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12552_ clknet_leaf_106_clk _01036_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11503_ _05703_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12483_ clknet_leaf_126_clk _00967_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11434_ _05295_ net559 _05657_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11365_ _05398_ rvsingle.dp.rf.rf\[14\]\[20\] _05618_ VGND VGND VPWR VPWR _05628_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_100_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_100_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13104_ clknet_leaf_51_clk _00562_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10316_ _04796_ net601 _05033_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__mux2_1
X_11296_ _05590_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__clkbuf_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ clknet_leaf_87_clk _00493_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10247_ _04996_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__clkbuf_1
X_10178_ _04929_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__buf_8
XFILLER_0_89_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12819_ clknet_leaf_35_clk _00277_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06340_ _01252_ _01254_ _01133_ _01262_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06271_ _01193_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08010_ rvsingle.dp.rf.rf\[19\]\[0\] _02929_ _02930_ VGND VGND VPWR VPWR _02931_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold603 rvsingle.dp.rf.rf\[29\]\[26\] VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold614 rvsingle.dp.rf.rf\[18\]\[18\] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold625 rvsingle.dp.rf.rf\[24\]\[19\] VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 rvsingle.dp.rf.rf\[5\]\[2\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 rvsingle.dp.rf.rf\[20\]\[14\] VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 rvsingle.dp.rf.rf\[16\]\[17\] VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09961_ _04779_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
Xhold669 rvsingle.dp.rf.rf\[9\]\[20\] VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08912_ _03778_ rvsingle.dp.rf.rf\[27\]\[25\] _03832_ VGND VGND VPWR VPWR _03833_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _04718_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__clkbuf_4
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _02211_ _02263_ _03763_ _02183_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__o31ai_2
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08774_ _01853_ _03689_ _03694_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__nand3_1
X_07725_ _01607_ rvsingle.dp.rf.rf\[20\]\[5\] VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__nor2_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07656_ _02534_ _02573_ _02576_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06607_ _01269_ rvsingle.dp.rf.rf\[16\]\[21\] VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07587_ rvsingle.dp.rf.rf\[17\]\[4\] _01267_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__or2b_1
X_09326_ _04239_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__nand2_1
X_06538_ rvsingle.dp.rf.rf\[1\]\[21\] _01441_ _01437_ VGND VGND VPWR VPWR _01459_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09257_ DataAdr[23] VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06469_ _01114_ _01388_ _01390_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08208_ _03128_ _02291_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09188_ _01134_ _04103_ _04107_ _01157_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08139_ Instr[27] _01084_ _01584_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_121_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11150_ _05510_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10101_ _04898_ net376 _04847_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__mux2_1
X_11081_ _05475_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__clkbuf_1
X_10032_ _04365_ _04837_ _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_98_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_149_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_149_clk sky130_fd_sc_hd__clkbuf_16
X_11983_ _05958_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10934_ _05393_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10865_ _05085_ _05350_ _05325_ net145 VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12604_ clknet_leaf_149_clk _00062_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10796_ _05307_ net517 _05298_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ clknet_leaf_15_clk _01019_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12466_ clknet_leaf_27_clk _00950_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11417_ _05645_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__buf_8
XFILLER_0_22_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12397_ clknet_leaf_43_clk _00881_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11348_ _05619_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11279_ _05207_ net438 _05580_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__mux2_1
X_13018_ clknet_leaf_12_clk _00476_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07510_ _02375_ Instr[26] VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08490_ _03409_ _03410_ _02329_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07441_ rvsingle.dp.rf.rf\[23\]\[7\] _01561_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__and2b_1
XFILLER_0_159_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07372_ _02274_ _02280_ _02284_ _02292_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09111_ _04017_ _04023_ _01378_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06323_ _01242_ _01244_ _01245_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__or3_4
XFILLER_0_33_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09042_ _01643_ rvsingle.dp.rf.rf\[4\]\[27\] VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__or2_1
X_06254_ Instr[5] _01063_ _01078_ _01067_ _01081_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_72_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold400 rvsingle.dp.rf.rf\[4\]\[14\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 rvsingle.dp.rf.rf\[21\]\[24\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
X_06185_ rvsingle.dp.rf.rf\[7\]\[30\] _01090_ _01108_ VGND VGND VPWR VPWR _01109_
+ sky130_fd_sc_hd__o21ai_1
Xhold422 rvsingle.dp.rf.rf\[10\]\[21\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold433 rvsingle.dp.rf.rf\[6\]\[8\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 rvsingle.dp.rf.rf\[29\]\[7\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 rvsingle.dp.rf.rf\[31\]\[10\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 rvsingle.dp.rf.rf\[8\]\[26\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 rvsingle.dp.rf.rf\[23\]\[25\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ _04765_ rvsingle.dp.rf.rf\[2\]\[5\] _04741_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__mux2_1
Xhold488 rvsingle.dp.rf.rf\[13\]\[13\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 rvsingle.dp.rf.rf\[21\]\[1\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _04618_ PC[31] VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__nand2_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _03397_ _03382_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__nand2_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _03676_ _03677_ _01111_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ rvsingle.dp.rf.rf\[3\]\[5\] _01606_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__or2b_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _01382_ rvsingle.dp.rf.rf\[16\]\[14\] VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__nor2_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _01721_ _02557_ _02559_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__nand3_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10650_ _04886_ net662 _05219_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09309_ _04224_ _03744_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10581_ _04898_ _05183_ _05146_ _05186_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12320_ _06111_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12251_ _06077_ net89 _05161_ _05832_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11202_ _05539_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12182_ _05004_ _05350_ _06052_ net177 VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__a2bb2o_1
X_11133_ _05385_ net533 _05499_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__mux2_1
X_11064_ _05330_ net374 _05460_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__mux2_1
X_10015_ _04824_ net687 _04791_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__mux2_1
X_11966_ _04781_ net751 _05949_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10917_ _05383_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__clkbuf_1
X_11897_ _04785_ net329 _05902_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10848_ _04802_ _05183_ _05336_ _05341_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10779_ _05297_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12518_ clknet_leaf_108_clk _01002_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12449_ clknet_leaf_141_clk _00933_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07990_ _01067_ _02909_ _02910_ _01173_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__nor4_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06941_ _01557_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__buf_8
XFILLER_0_158_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09660_ _01171_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__clkbuf_4
X_06872_ _01126_ rvsingle.dp.rf.rf\[18\]\[23\] _01105_ _01792_ VGND VGND VPWR VPWR
+ _01793_ sky130_fd_sc_hd__o211a_1
X_08611_ rvsingle.dp.rf.rf\[1\]\[12\] _01561_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__and2b_1
X_09591_ _04429_ PC[6] _04421_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__and3_1
X_08542_ _01349_ rvsingle.dp.rf.rf\[28\]\[13\] VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08473_ rvsingle.dp.rf.rf\[17\]\[9\] _01827_ _01308_ _03393_ VGND VGND VPWR VPWR
+ _03394_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_65_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07424_ _02336_ _02339_ _01156_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07355_ _01725_ rvsingle.dp.rf.rf\[8\]\[7\] _01299_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06306_ _01172_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07286_ rvsingle.dp.rf.rf\[8\]\[16\] rvsingle.dp.rf.rf\[9\]\[16\] rvsingle.dp.rf.rf\[10\]\[16\]
+ rvsingle.dp.rf.rf\[11\]\[16\] _01707_ _01244_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09025_ rvsingle.dp.rf.rf\[21\]\[27\] _01089_ _01093_ _03944_ VGND VGND VPWR VPWR
+ _03945_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06237_ rvsingle.dp.rf.rf\[28\]\[30\] rvsingle.dp.rf.rf\[29\]\[30\] _01128_ VGND
+ VGND VPWR VPWR _01161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold230 rvsingle.dp.rf.rf\[6\]\[22\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 rvsingle.dp.rf.rf\[4\]\[19\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ _01091_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__buf_8
XFILLER_0_130_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold252 rvsingle.dp.rf.rf\[4\]\[28\] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 rvsingle.dp.rf.rf\[12\]\[30\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 rvsingle.dp.rf.rf\[27\]\[24\] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 rvsingle.dp.rf.rf\[19\]\[29\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 rvsingle.dp.rf.rf\[1\]\[26\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09927_ _04750_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__buf_4
X_09858_ _04685_ _04686_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__nand3_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _03696_ _01481_ _02505_ _03673_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__nand4_2
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _04398_ _04616_ _04624_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[23\] sky130_fd_sc_hd__o21ai_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _01215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11820_ _05740_ net270 _05863_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__mux2_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _01426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 _01493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _01520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _01595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _05839_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_158 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_169 _01699_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
X_10702_ _05254_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _05534_ rvsingle.dp.rf.rf\[10\]\[5\] _05795_ VGND VGND VPWR VPWR _05800_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _04834_ net507 _05205_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13352_ clknet_leaf_80_clk rvsingle.dp.PCNext\[29\] _00029_ VGND VGND VPWR VPWR PC[29]
+ sky130_fd_sc_hd__dfrtp_4
X_10564_ _05167_ _05177_ _05155_ net186 VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12303_ _06102_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13283_ clknet_leaf_125_clk _00741_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10495_ _05135_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12234_ reset VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12165_ _06053_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
X_11116_ _05492_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__clkbuf_1
X_12096_ _06017_ _05060_ _04924_ _06010_ net33 VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a32o_1
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11047_ _05145_ _05457_ net108 VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__a21oi_1
X_12998_ clknet_leaf_115_clk _00456_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11949_ _05724_ rvsingle.dp.rf.rf\[4\]\[1\] _05940_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_71_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07140_ rvsingle.dp.rf.rf\[11\]\[18\] _01540_ _02060_ VGND VGND VPWR VPWR _02061_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07071_ _01656_ rvsingle.dp.rf.rf\[14\]\[19\] _01605_ VGND VGND VPWR VPWR _01992_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07973_ rvsingle.dp.rf.rf\[26\]\[0\] _01562_ _02320_ _02893_ VGND VGND VPWR VPWR
+ _02894_ sky130_fd_sc_hd__o211ai_1
X_09712_ PC[16] _04543_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__nor2_1
X_06924_ rvsingle.dp.rf.rf\[13\]\[22\] _01088_ _01668_ VGND VGND VPWR VPWR _01845_
+ sky130_fd_sc_hd__o21ai_1
X_09643_ _04140_ MemWrite _01090_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__o21ai_1
X_06855_ _01744_ rvsingle.dp.rf.rf\[26\]\[23\] _01648_ _01775_ VGND VGND VPWR VPWR
+ _01776_ sky130_fd_sc_hd__o211a_1
X_09574_ _04367_ _04420_ _04421_ _04428_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[4\]
+ sky130_fd_sc_hd__o2bb2ai_1
X_06786_ _01419_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__buf_6
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _01642_ rvsingle.dp.rf.rf\[4\]\[13\] VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08456_ rvsingle.dp.rf.rf\[5\]\[9\] _01827_ _01308_ _03376_ VGND VGND VPWR VPWR _03377_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_136_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07407_ rvsingle.dp.rf.rf\[9\]\[7\] _01136_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08387_ _03305_ _01716_ _01460_ _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07338_ Instr[4] VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07269_ _02186_ _02188_ _01208_ _02189_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09008_ _01302_ _03927_ _01230_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10280_ _05014_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__clkbuf_1
X_12921_ clknet_leaf_8_clk _00379_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ clknet_leaf_21_clk _00310_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _05721_ _05860_ _05861_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__a21oi_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ clknet_leaf_66_clk _00241_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ _05639_ net452 _05817_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__mux2_1
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11665_ _04904_ _05766_ _05457_ _05789_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__a31o_1
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13404_ clknet_leaf_147_clk _00832_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10616_ _04794_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__buf_2
XFILLER_0_92_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11596_ _04863_ _04973_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13335_ clknet_leaf_75_clk rvsingle.dp.PCNext\[12\] _00012_ VGND VGND VPWR VPWR PC[12]
+ sky130_fd_sc_hd__dfrtp_4
X_10547_ _05167_ _05168_ _05155_ net114 VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_45_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13266_ clknet_leaf_67_clk _00724_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10478_ _05102_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__buf_8
X_12217_ _06068_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__inv_2
X_13197_ clknet_leaf_90_clk _00655_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12148_ _04720_ _04725_ _04967_ _04968_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__and4_2
X_12079_ _05316_ _05099_ net147 VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06640_ _01135_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__buf_6
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06571_ _01135_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_16
X_08310_ _03141_ net821 _03221_ _03227_ _03230_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__o2111ai_4
X_09290_ _04203_ _04204_ _04137_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08241_ rvsingle.dp.rf.rf\[4\]\[10\] rvsingle.dp.rf.rf\[5\]\[10\] rvsingle.dp.rf.rf\[6\]\[10\]
+ rvsingle.dp.rf.rf\[7\]\[10\] _01416_ _01708_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__mux4_1
XANTENNA_14 DataAdr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 Instr[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_36 Instr[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 ReadData[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ _02005_ rvsingle.dp.rf.rf\[0\]\[11\] _01519_ VGND VGND VPWR VPWR _03093_
+ sky130_fd_sc_hd__o21bai_1
XANTENNA_69 ReadData[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07123_ _01630_ rvsingle.dp.rf.rf\[4\]\[18\] VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_928 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07054_ rvsingle.dp.rf.rf\[25\]\[19\] _01862_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07956_ rvsingle.dp.rf.rf\[8\]\[0\] _01619_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__nor2_1
X_06907_ _01190_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__buf_6
X_07887_ _02805_ _02273_ _02807_ _01217_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06838_ _01667_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__buf_4
X_09626_ PC[8] _04456_ PC[9] VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09557_ _04398_ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__nand2_1
X_06769_ _01190_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__buf_4
XFILLER_0_167_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
X_08508_ _03417_ _03428_ _01145_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__nand3_4
X_09488_ _01154_ _01641_ _01683_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__and3_2
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08439_ rvsingle.dp.rf.rf\[23\]\[9\] _01492_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__or2b_1
XFILLER_0_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11450_ _05674_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10401_ _05064_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__buf_8
XFILLER_0_135_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11381_ _05636_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13120_ clknet_leaf_138_clk _00578_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10332_ _04840_ net718 _05033_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13051_ clknet_leaf_131_clk _00509_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10263_ _04981_ _04839_ _04982_ _04983_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__and4b_2
XFILLER_0_103_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12002_ _05713_ net225 _05960_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__mux2_1
X_10194_ _04960_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12904_ clknet_leaf_105_clk _00362_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12835_ clknet_leaf_127_clk _00293_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12766_ clknet_leaf_150_clk _00224_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11717_ _05818_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ clknet_leaf_23_clk _00155_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11648_ net65 _05778_ _05754_ _05457_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11579_ _05344_ net690 _05729_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold807 rvsingle.dp.rf.rf\[20\]\[4\] VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_124_clk _00776_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold818 rvsingle.dp.rf.rf\[25\]\[13\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13249_ clknet_leaf_128_clk _00707_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07810_ _02337_ _02727_ _02728_ _01599_ _02730_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__o311ai_1
X_08790_ _01721_ _03708_ _03710_ _01446_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__a31oi_1
X_07741_ _01150_ _01139_ _02657_ _02633_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__o211ai_4
X_07672_ _02582_ _02586_ _02590_ _02592_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__o22ai_4
X_09411_ _02211_ _04322_ _04247_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__a21o_1
X_06623_ _01095_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
X_09342_ _03565_ _03567_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__nand2_1
X_06554_ _01192_ rvsingle.dp.rf.rf\[12\]\[21\] VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09273_ _04187_ _04189_ VGND VGND VPWR VPWR DataAdr[30] sky130_fd_sc_hd__nand2_8
X_06485_ _01066_ _01075_ _01405_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__or3b_2
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08224_ _01422_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08155_ _01743_ rvsingle.dp.rf.rf\[24\]\[11\] _01519_ VGND VGND VPWR VPWR _03076_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_16_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07106_ _02021_ _02026_ _01526_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__nand3_1
XFILLER_0_43_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08086_ _03004_ _03006_ _01502_ _01115_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07037_ _01218_ _01949_ _01957_ _01316_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_140_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08988_ _03880_ _03881_ _03907_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__o21ai_2
X_07939_ _01065_ _01074_ _01870_ _02849_ _02798_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__o221a_1
X_10950_ _05300_ rvsingle.dp.rf.rf\[18\]\[22\] _05401_ VGND VGND VPWR VPWR _05403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09609_ _04451_ _04453_ _04460_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[7\] sky130_fd_sc_hd__o21ai_1
X_10881_ _05359_ net641 _05319_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12620_ clknet_leaf_50_clk _00078_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12551_ clknet_leaf_127_clk _01035_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11502_ _05439_ net628 _05695_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12482_ clknet_leaf_128_clk _00966_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11433_ _05665_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11364_ _05627_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10315_ _05034_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__clkbuf_1
X_13103_ clknet_leaf_58_clk _00561_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11295_ _05398_ net788 _05580_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ clknet_leaf_93_clk _00492_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10246_ _04802_ net763 _04989_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10177_ _04951_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12818_ clknet_leaf_47_clk _00276_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12749_ clknet_leaf_43_clk _00207_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06270_ _01192_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__buf_4
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold604 rvsingle.dp.rf.rf\[14\]\[14\] VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold615 rvsingle.dp.rf.rf\[2\]\[19\] VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold626 rvsingle.dp.rf.rf\[24\]\[20\] VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 rvsingle.dp.rf.rf\[31\]\[25\] VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 rvsingle.dp.rf.rf\[2\]\[13\] VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold659 rvsingle.dp.rf.rf\[25\]\[2\] VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _04778_ net676 _04741_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_6_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08911_ _01848_ rvsingle.dp.rf.rf\[26\]\[25\] _01648_ VGND VGND VPWR VPWR _03832_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09891_ PC[0] _04426_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__o21ai_4
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _01581_ _02262_ _01837_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__a21oi_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _01660_ _03690_ _03691_ _02410_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__o311ai_1
X_07724_ rvsingle.dp.rf.rf\[21\]\[5\] VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ _02469_ _02574_ _02534_ _02575_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06606_ _01522_ _01112_ _01525_ _01526_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_94_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07586_ rvsingle.dp.rf.rf\[19\]\[4\] _02481_ _01552_ VGND VGND VPWR VPWR _02507_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09325_ _04240_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06537_ _01193_ rvsingle.dp.rf.rf\[0\]\[21\] VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09256_ _01804_ _04144_ _04174_ VGND VGND VPWR VPWR DataAdr[23] sky130_fd_sc_hd__o21ai_4
X_06468_ _01133_ _01389_ _01157_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08207_ rvsingle.dp.rf.rf\[21\]\[11\] _02303_ _01308_ _03127_ VGND VGND VPWR VPWR
+ _03128_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_145_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09187_ _01120_ _04104_ _04106_ _01114_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06399_ rvsingle.dp.rf.rf\[14\]\[29\] rvsingle.dp.rf.rf\[15\]\[29\] _01195_ VGND
+ VGND VPWR VPWR _01321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08138_ _01592_ _02346_ _02371_ _01178_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__a31o_1
XFILLER_0_160_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08069_ _01695_ rvsingle.dp.rf.rf\[30\]\[1\] VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__nor2_1
X_10100_ _04897_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11080_ _05291_ rvsingle.dp.rf.rf\[17\]\[16\] _05469_ VGND VGND VPWR VPWR _05475_
+ sky130_fd_sc_hd__mux2_1
X_10031_ _04505_ _04506_ _04595_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__and3_1
X_11982_ _04823_ net321 _05949_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10933_ _05212_ rvsingle.dp.rf.rf\[18\]\[15\] _05387_ VGND VGND VPWR VPWR _05393_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10864_ _04846_ _05316_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12603_ clknet_leaf_142_clk _00061_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10795_ _04885_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__buf_2
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_783 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ clknet_leaf_35_clk _01018_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12465_ clknet_leaf_48_clk _00949_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11416_ _05656_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__clkbuf_1
X_12396_ clknet_leaf_50_clk _00880_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11347_ _05334_ net468 _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11278_ _05581_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13017_ clknet_leaf_10_clk _00475_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10229_ _04981_ _04764_ _04982_ _04983_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__and4b_1
Xhold1 rvsingle.dp.rf.rf\[9\]\[0\] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07440_ _01675_ rvsingle.dp.rf.rf\[22\]\[7\] _01654_ VGND VGND VPWR VPWR _02361_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07371_ _02287_ _02290_ _02291_ _01446_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__a31o_1
X_09110_ _01133_ _04024_ _04029_ _01117_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_72_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06322_ Instr[17] _01215_ Instr[19] VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__or3_2
XFILLER_0_128_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09041_ _02236_ _03958_ _03960_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06253_ _01172_ _01076_ _01175_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold401 rvsingle.dp.rf.rf\[30\]\[24\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06184_ _01100_ rvsingle.dp.rf.rf\[6\]\[30\] _01107_ VGND VGND VPWR VPWR _01108_
+ sky130_fd_sc_hd__o21a_1
Xhold412 rvsingle.dp.rf.rf\[10\]\[18\] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold423 rvsingle.dp.rf.rf\[21\]\[12\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 rvsingle.dp.rf.rf\[28\]\[11\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 rvsingle.dp.rf.rf\[24\]\[4\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold456 rvsingle.dp.rf.rf\[26\]\[22\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold467 rvsingle.dp.rf.rf\[12\]\[9\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 rvsingle.dp.rf.rf\[9\]\[17\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _04764_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__buf_2
Xhold489 rvsingle.dp.rf.rf\[1\]\[10\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _04618_ PC[31] VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__or2_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ net821 _03141_ _03227_ _03221_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__o211a_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ rvsingle.dp.rf.rf\[9\]\[15\] _01613_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__or2b_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ rvsingle.dp.rf.rf\[1\]\[5\] _02627_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _03602_ _03607_ _02527_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__nand3_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ rvsingle.dp.rf.rf\[27\]\[4\] _01901_ _02558_ VGND VGND VPWR VPWR _02559_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07569_ _01493_ rvsingle.dp.rf.rf\[6\]\[4\] _01552_ _02489_ VGND VGND VPWR VPWR _02490_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09308_ _04220_ _04223_ _03650_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10580_ _05085_ _05149_ net535 VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09239_ _04154_ _04157_ _03062_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_161_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12250_ _06077_ net129 _05466_ _05832_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11201_ _05428_ net404 _05528_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12181_ _04840_ _05766_ _05336_ _06057_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11132_ _05490_ net123 _05116_ _05501_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__a22o_1
X_11063_ _05463_ net135 _05161_ _05464_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__a22o_1
X_10014_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__buf_2
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11965_ _05939_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__buf_6
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10916_ _05330_ net555 _05373_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11896_ _05911_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10847_ _05337_ _05338_ _05339_ _05084_ net195 VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__o41a_1
XFILLER_0_128_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10778_ _04840_ net794 _05285_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12517_ clknet_leaf_115_clk _01001_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12448_ clknet_leaf_120_clk _00932_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12379_ clknet_leaf_136_clk _00863_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06940_ _01860_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06871_ rvsingle.dp.rf.rf\[19\]\[23\] _01753_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__or2b_1
XFILLER_0_94_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08610_ _01630_ rvsingle.dp.rf.rf\[0\]\[12\] VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__nor2_1
X_09590_ _04441_ _04442_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__nor2_1
X_08541_ _01440_ rvsingle.dp.rf.rf\[31\]\[13\] _02162_ _03461_ VGND VGND VPWR VPWR
+ _03462_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08472_ _02163_ rvsingle.dp.rf.rf\[16\]\[9\] VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07423_ _01552_ _02340_ _02341_ _01111_ _02343_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_147_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07354_ _01294_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06305_ _01210_ _01227_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07285_ rvsingle.dp.rf.rf\[12\]\[16\] rvsingle.dp.rf.rf\[13\]\[16\] rvsingle.dp.rf.rf\[14\]\[16\]
+ rvsingle.dp.rf.rf\[15\]\[16\] _01336_ _01200_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09024_ _01643_ rvsingle.dp.rf.rf\[20\]\[27\] VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__or2_1
X_06236_ _01158_ _01159_ _01114_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold220 rvsingle.dp.rf.rf\[16\]\[22\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06167_ Instr[21] VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__inv_2
Xhold231 rvsingle.dp.rf.rf\[5\]\[11\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 rvsingle.dp.rf.rf\[8\]\[23\] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 rvsingle.dp.rf.rf\[12\]\[2\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold264 rvsingle.dp.rf.rf\[5\]\[28\] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 rvsingle.dp.rf.rf\[4\]\[4\] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold286 rvsingle.dp.rf.rf\[28\]\[28\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 rvsingle.dp.rf.rf\[26\]\[28\] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__buf_4
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _04617_ PC[29] VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__nand2_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _03699_ _03727_ _03728_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__nand3_2
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _04366_ _04622_ _04623_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__nand3_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _01218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08739_ _03656_ _03657_ _03659_ _02488_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__o211ai_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _01426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _01499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _01531_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _01605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _05728_ net799 _05837_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__mux2_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _01675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _04828_ net521 _05246_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__mux2_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _05799_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10632_ _05216_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10563_ _04846_ _05144_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__nand2_1
X_13351_ clknet_leaf_79_clk rvsingle.dp.PCNext\[28\] _00028_ VGND VGND VPWR VPWR PC[28]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12302_ _04754_ net610 _06099_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__mux2_1
X_13282_ clknet_leaf_119_clk _00740_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10494_ _04877_ net462 _05126_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12233_ reset VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12164_ _05740_ net511 _06049_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11115_ _05322_ net572 _05490_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__mux2_1
X_12095_ _04773_ _04726_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__and2_1
X_11046_ _05367_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12997_ clknet_leaf_108_clk _00455_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11948_ _05939_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__buf_6
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11879_ _05724_ rvsingle.dp.rf.rf\[6\]\[1\] _05902_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07070_ rvsingle.dp.rf.rf\[15\]\[19\] VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07972_ rvsingle.dp.rf.rf\[27\]\[0\] _01561_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09711_ PC[14] PC[15] PC[16] _04522_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__and4_1
X_06923_ _01098_ rvsingle.dp.rf.rf\[12\]\[22\] VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__nor2_1
X_09642_ _04367_ _04480_ _04490_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[10\] sky130_fd_sc_hd__o21ai_1
X_06854_ rvsingle.dp.rf.rf\[27\]\[23\] _01753_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__or2b_1
XFILLER_0_117_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06785_ _01625_ _01329_ _01199_ _01705_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__a211o_1
X_09573_ _04422_ _04423_ _04424_ _04427_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_117_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _01520_ _03441_ _03442_ _01564_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08455_ _02163_ rvsingle.dp.rf.rf\[4\]\[9\] VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07406_ _01148_ rvsingle.dp.rf.rf\[8\]\[7\] VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08386_ _02929_ rvsingle.dp.rf.rf\[23\]\[8\] _03306_ VGND VGND VPWR VPWR _03307_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07337_ _02257_ _01482_ _01837_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07268_ rvsingle.dp.rf.rf\[20\]\[16\] rvsingle.dp.rf.rf\[21\]\[16\] rvsingle.dp.rf.rf\[22\]\[16\]
+ rvsingle.dp.rf.rf\[23\]\[16\] _01432_ _01434_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09007_ rvsingle.dp.rf.rf\[10\]\[27\] rvsingle.dp.rf.rf\[11\]\[27\] _01242_ VGND
+ VGND VPWR VPWR _03927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06219_ _01114_ _01123_ _01142_ _01118_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07199_ _01848_ rvsingle.dp.rf.rf\[20\]\[17\] VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09909_ PC[1] _04425_ _04731_ _04734_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__o22a_4
X_12920_ clknet_leaf_32_clk _00378_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ clknet_leaf_35_clk _00309_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11802_ net120 _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__nor2_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12782_ clknet_leaf_68_clk _00240_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11733_ _05826_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__clkbuf_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _04976_ _05417_ _05371_ net518 VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__o31a_1
XFILLER_0_138_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13403_ clknet_leaf_142_clk _00831_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10615_ _05206_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__clkbuf_1
X_11595_ _05758_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13334_ clknet_leaf_75_clk rvsingle.dp.PCNext\[11\] _00011_ VGND VGND VPWR VPWR PC[11]
+ sky130_fd_sc_hd__dfrtp_4
X_10546_ _04802_ _05145_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13265_ clknet_leaf_55_clk _00723_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10477_ _05125_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12216_ _06068_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__inv_2
X_13196_ clknet_leaf_93_clk _00654_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12147_ _06043_ _06007_ _06044_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__o21ai_1
X_12078_ _04721_ _04726_ _04924_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__and3_1
X_11029_ _05447_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06570_ _01490_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08240_ _02302_ _03155_ _03160_ _02438_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_28_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 DataAdr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 Instr[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 Instr[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08171_ _01552_ _03088_ _03089_ _02323_ _03091_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__o311a_1
XFILLER_0_133_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_59 ReadData[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07122_ rvsingle.dp.rf.rf\[7\]\[18\] _01861_ _01260_ VGND VGND VPWR VPWR _02043_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07053_ _01656_ rvsingle.dp.rf.rf\[24\]\[19\] VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07955_ rvsingle.dp.rf.rf\[9\]\[0\] VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__inv_2
X_06906_ _01294_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__clkbuf_8
X_07886_ rvsingle.dp.rf.rf\[15\]\[2\] _02275_ _02806_ VGND VGND VPWR VPWR _02807_
+ sky130_fd_sc_hd__o21ai_1
X_09625_ PC[8] PC[9] _04456_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__and3_2
X_06837_ rvsingle.dp.rf.rf\[7\]\[23\] VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09556_ _04409_ _04411_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__xor2_1
X_06768_ _01307_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__buf_6
XFILLER_0_167_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08507_ _03420_ _03422_ _02364_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_78_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09487_ _04384_ VGND VGND VPWR VPWR WriteData[21] sky130_fd_sc_hd__clkbuf_4
X_06699_ _01530_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__buf_6
XFILLER_0_163_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08438_ rvsingle.dp.rf.rf\[21\]\[9\] _01125_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08369_ rvsingle.dp.rf.rf\[12\]\[8\] rvsingle.dp.rf.rf\[13\]\[8\] rvsingle.dp.rf.rf\[14\]\[8\]
+ rvsingle.dp.rf.rf\[15\]\[8\] _01241_ _01953_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10400_ _05000_ _05068_ _05069_ _05065_ net10 VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11380_ _05307_ net728 _05629_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10331_ _05042_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10262_ _05004_ _05005_ _04978_ net156 VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__a2bb2o_1
X_13050_ clknet_leaf_12_clk _00508_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12001_ _05967_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__clkbuf_1
X_10193_ _04892_ net286 _04952_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12903_ clknet_leaf_98_clk _00361_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12834_ clknet_leaf_129_clk _00292_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ clknet_leaf_143_clk _00223_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _04845_ net422 _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__mux2_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ clknet_leaf_19_clk _00154_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11647_ _05371_ _05753_ _05779_ net133 VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_126_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11578_ _05167_ _05749_ _05731_ net104 VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_52_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold808 rvsingle.dp.rf.rf\[7\]\[1\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13317_ clknet_leaf_126_clk _00775_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10529_ _05113_ _05114_ _05115_ _05061_ _04764_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__o311a_1
X_13248_ clknet_leaf_134_clk _00706_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13179_ clknet_leaf_18_clk _00637_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_07740_ _02469_ _02608_ _02659_ _02660_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07671_ _01721_ _02591_ _02438_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__o21ai_1
X_09410_ _02257_ _01085_ _01837_ _03142_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__a211o_1
X_06622_ _01542_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06553_ _01441_ rvsingle.dp.rf.rf\[15\]\[21\] _01434_ _01473_ VGND VGND VPWR VPWR
+ _01474_ sky130_fd_sc_hd__o211a_1
X_09341_ _03565_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06484_ _01085_ WriteData[28] _01180_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__a21o_1
X_09272_ _04121_ _04188_ _04122_ _01186_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__or4b_4
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08223_ rvsingle.dp.rf.rf\[20\]\[10\] rvsingle.dp.rf.rf\[21\]\[10\] rvsingle.dp.rf.rf\[22\]\[10\]
+ rvsingle.dp.rf.rf\[23\]\[10\] _02176_ _01696_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08154_ _01156_ _03069_ _03074_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__nand3_1
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07105_ _02022_ _02023_ _01112_ _02025_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08085_ _01797_ rvsingle.dp.rf.rf\[6\]\[1\] _01647_ _03005_ VGND VGND VPWR VPWR _03006_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_3_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07036_ _01208_ _01950_ _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08987_ _01351_ _01203_ _03892_ _03906_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__o211ai_4
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07938_ _01316_ _02814_ _02825_ _01452_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__a31o_1
X_07869_ _01490_ _02786_ _02787_ _02329_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09608_ _04454_ _04455_ _04458_ _04459_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_168_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10880_ _04891_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09539_ _04138_ _04132_ VGND VGND VPWR VPWR DataAdr[31] sky130_fd_sc_hd__nand2_8
XFILLER_0_78_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12550_ clknet_leaf_108_clk _01034_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11501_ _05702_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12481_ clknet_leaf_140_clk _00965_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11432_ _05439_ net713 _05657_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11363_ _05295_ net725 _05618_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ clknet_leaf_55_clk _00560_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10314_ _04790_ net353 _05033_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__mux2_1
X_11294_ _05589_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ clknet_leaf_90_clk _00491_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10245_ _04995_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__clkbuf_1
X_10176_ _04840_ net273 _04941_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12817_ clknet_leaf_48_clk _00275_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12748_ clknet_leaf_50_clk _00206_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12679_ clknet_leaf_104_clk _00137_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold605 rvsingle.dp.rf.rf\[2\]\[21\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold616 rvsingle.dp.rf.rf\[25\]\[29\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 rvsingle.dp.rf.rf\[12\]\[6\] VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 rvsingle.dp.rf.rf\[1\]\[2\] VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 rvsingle.dp.rf.rf\[7\]\[8\] VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
X_08910_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _01169_ _01170_ _02259_ _04714_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__o32ai_4
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _03142_ _03761_ _02151_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _02030_ rvsingle.dp.rf.rf\[6\]\[15\] _02337_ _03692_ VGND VGND VPWR VPWR
+ _03693_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_109_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07723_ _02638_ _02643_ _02491_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__nand3_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07654_ _02473_ _02318_ _01537_ _02571_ _02530_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__o221a_1
X_06605_ _01115_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__buf_6
XFILLER_0_76_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07585_ _01518_ rvsingle.dp.rf.rf\[18\]\[4\] VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09324_ _03909_ _03908_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__nand2_1
X_06536_ rvsingle.dp.rf.rf\[4\]\[21\] rvsingle.dp.rf.rf\[5\]\[21\] rvsingle.dp.rf.rf\[6\]\[21\]
+ rvsingle.dp.rf.rf\[7\]\[21\] _01329_ _01456_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__mux4_1
XFILLER_0_168_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09255_ _01840_ _04170_ _04173_ _04137_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__o211ai_2
X_06467_ rvsingle.dp.rf.rf\[20\]\[28\] rvsingle.dp.rf.rf\[21\]\[28\] rvsingle.dp.rf.rf\[22\]\[28\]
+ rvsingle.dp.rf.rf\[23\]\[28\] _01138_ _01106_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08206_ _01191_ rvsingle.dp.rf.rf\[20\]\[11\] VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06398_ rvsingle.dp.rf.rf\[13\]\[29\] _01298_ _01311_ _01319_ VGND VGND VPWR VPWR
+ _01320_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09186_ rvsingle.dp.rf.rf\[1\]\[31\] _01090_ _01094_ _04105_ VGND VGND VPWR VPWR
+ _04106_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08137_ _03056_ _02667_ _03057_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08068_ rvsingle.dp.rf.rf\[24\]\[1\] rvsingle.dp.rf.rf\[25\]\[1\] rvsingle.dp.rf.rf\[26\]\[1\]
+ rvsingle.dp.rf.rf\[27\]\[1\] _01903_ _01470_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07019_ _01939_ _01309_ _01207_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10030_ _02908_ DataAdr[20] _04836_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11981_ _05957_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__clkbuf_1
X_10932_ _05392_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10863_ _04840_ _05183_ _05336_ _05349_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12602_ clknet_leaf_3_clk _00060_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10794_ _05306_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__clkbuf_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12533_ clknet_leaf_36_clk _01017_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12464_ clknet_leaf_70_clk _00948_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11415_ _05385_ rvsingle.dp.rf.rf\[13\]\[10\] _05646_ VGND VGND VPWR VPWR _05656_
+ sky130_fd_sc_hd__mux2_1
X_12395_ clknet_leaf_87_clk _00879_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11346_ _05606_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__buf_8
XFILLER_0_10_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11277_ _05334_ net717 _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13016_ clknet_leaf_23_clk _00474_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10228_ _04986_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 rvsingle.dp.rf.rf\[25\]\[5\] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _04942_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07370_ _01172_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06321_ _01243_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__buf_6
XFILLER_0_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09040_ rvsingle.dp.rf.rf\[3\]\[27\] _03778_ _03959_ VGND VGND VPWR VPWR _03960_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06252_ _01173_ _01174_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__nor2_4
XFILLER_0_60_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06183_ _01106_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold402 rvsingle.dp.rf.rf\[22\]\[30\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold413 rvsingle.dp.rf.rf\[20\]\[24\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 rvsingle.dp.rf.rf\[20\]\[23\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold435 rvsingle.dp.rf.rf\[5\]\[17\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 rvsingle.dp.rf.rf\[26\]\[29\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold457 rvsingle.dp.rf.rf\[26\]\[14\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 rvsingle.dp.rf.rf\[14\]\[11\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09942_ _04426_ _04762_ _04763_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__a21o_4
Xhold479 rvsingle.dp.rf.rf\[22\]\[9\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _04618_ PC[30] VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__and2_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _03737_ _03740_ _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__nand3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _01561_ rvsingle.dp.rf.rf\[8\]\[15\] _01489_ VGND VGND VPWR VPWR _03676_
+ sky130_fd_sc_hd__o21ba_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _01135_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__clkbuf_8
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _01605_ _03603_ _03604_ _02351_ _03606_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _01903_ rvsingle.dp.rf.rf\[26\]\[4\] _01243_ VGND VGND VPWR VPWR _02558_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07568_ rvsingle.dp.rf.rf\[7\]\[4\] _01618_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09307_ _03572_ _03755_ _04222_ _03737_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06519_ _01294_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__clkbuf_8
X_07499_ _01097_ rvsingle.dp.rf.rf\[4\]\[6\] VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09238_ _03056_ _02667_ _03057_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09169_ rvsingle.dp.rf.rf\[30\]\[31\] rvsingle.dp.rf.rf\[31\]\[31\] _02212_ VGND
+ VGND VPWR VPWR _04089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11200_ _05538_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__clkbuf_1
X_12180_ _05337_ _05338_ _05339_ _05003_ net192 VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__o41a_1
XFILLER_0_102_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11131_ _05367_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__buf_4
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11062_ net54 _05460_ _05466_ _05464_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__a22o_1
X_10013_ _04426_ _04821_ _04822_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__a21o_4
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11964_ _05948_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10915_ _05382_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__clkbuf_1
X_11895_ _05428_ net643 _05902_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10846_ _04796_ _05183_ _05336_ _05340_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10777_ _05296_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12516_ clknet_leaf_108_clk _01000_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12447_ clknet_leaf_13_clk _00931_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12378_ clknet_leaf_14_clk _00862_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11329_ _05609_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06870_ _01789_ _01790_ _01768_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08540_ _02163_ rvsingle.dp.rf.rf\[30\]\[13\] VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08471_ _01695_ rvsingle.dp.rf.rf\[18\]\[9\] _01433_ VGND VGND VPWR VPWR _03392_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07422_ _01658_ rvsingle.dp.rf.rf\[6\]\[7\] _01654_ _02342_ VGND VGND VPWR VPWR _02343_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07353_ _02267_ _02269_ _02270_ _02272_ _02273_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__o221a_2
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06304_ rvsingle.dp.rf.rf\[20\]\[30\] rvsingle.dp.rf.rf\[21\]\[30\] rvsingle.dp.rf.rf\[22\]\[30\]
+ rvsingle.dp.rf.rf\[23\]\[30\] _01225_ _01226_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07284_ _02191_ _02199_ _02204_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09023_ _03940_ _01093_ _01113_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_72_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06235_ rvsingle.dp.rf.rf\[20\]\[30\] rvsingle.dp.rf.rf\[21\]\[30\] rvsingle.dp.rf.rf\[22\]\[30\]
+ rvsingle.dp.rf.rf\[23\]\[30\] _01128_ _01107_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold210 rvsingle.dp.rf.rf\[1\]\[6\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 rvsingle.dp.rf.rf\[30\]\[28\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
X_06166_ _01089_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__buf_4
Xhold232 rvsingle.dp.rf.rf\[5\]\[16\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 rvsingle.dp.rf.rf\[4\]\[30\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 rvsingle.dp.rf.rf\[9\]\[24\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold265 rvsingle.dp.rf.rf\[0\]\[17\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold276 rvsingle.dp.rf.rf\[5\]\[29\] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 rvsingle.dp.rf.rf\[10\]\[29\] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold298 rvsingle.dp.rf.rf\[23\]\[1\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _01080_ _04121_ _01078_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__and3_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _04617_ PC[29] VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__or2_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _01960_ _02102_ _01961_ _03697_ _01580_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__o221ai_4
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _04607_ _04621_ _04619_ _04620_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__o211ai_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06999_ rvsingle.dp.rf.rf\[0\]\[22\] rvsingle.dp.rf.rf\[1\]\[22\] rvsingle.dp.rf.rf\[2\]\[22\]
+ rvsingle.dp.rf.rf\[3\]\[22\] _01432_ _01434_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__mux4_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _01878_ rvsingle.dp.rf.rf\[20\]\[15\] _03658_ _02395_ VGND VGND VPWR VPWR
+ _03659_ sky130_fd_sc_hd__o211ai_1
XANTENNA_105 _01247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _01427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _01499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _01545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_149 _01605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _01711_ _03589_ _01699_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__o21ai_2
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _05253_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _05377_ net598 _05795_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10631_ _04828_ net558 _05205_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13350_ clknet_leaf_79_clk rvsingle.dp.PCNext\[27\] _00027_ VGND VGND VPWR VPWR PC[27]
+ sky130_fd_sc_hd__dfrtp_4
X_10562_ _05176_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12301_ _06101_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13281_ clknet_leaf_131_clk _00739_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10493_ _05134_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12232_ _06069_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12163_ net19 _06052_ _06017_ _04985_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11114_ _05491_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__clkbuf_1
X_12094_ _06016_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__clkbuf_1
X_11045_ _04721_ _05058_ _05367_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__and3_2
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12996_ clknet_leaf_109_clk _00454_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11947_ _04737_ _04739_ _04976_ _05835_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__or4_2
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__buf_6
XFILLER_0_156_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10829_ _04774_ net383 _05320_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07971_ rvsingle.dp.rf.rf\[25\]\[0\] _01796_ _02891_ VGND VGND VPWR VPWR _02892_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09710_ _04547_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__xnor2_1
X_06922_ rvsingle.dp.rf.rf\[15\]\[22\] _01842_ _01612_ VGND VGND VPWR VPWR _01843_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09641_ _04366_ _04487_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__nand3_1
X_06853_ _01593_ _01757_ _01773_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__nand3_2
X_09572_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__clkbuf_4
X_06784_ _01420_ rvsingle.dp.rf.rf\[4\]\[20\] VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08523_ _01642_ rvsingle.dp.rf.rf\[2\]\[13\] _01596_ _03443_ VGND VGND VPWR VPWR
+ _03444_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_148_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08454_ rvsingle.dp.rf.rf\[0\]\[9\] rvsingle.dp.rf.rf\[1\]\[9\] rvsingle.dp.rf.rf\[2\]\[9\]
+ rvsingle.dp.rf.rf\[3\]\[9\] _02176_ _02162_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07405_ _02320_ _02321_ _02322_ _02323_ _02325_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__o311ai_4
X_08385_ _01240_ rvsingle.dp.rf.rf\[22\]\[8\] _01454_ VGND VGND VPWR VPWR _03306_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07336_ _01962_ _02212_ _02234_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_46_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07267_ _02187_ _01717_ _01703_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09006_ _03924_ _01330_ _01451_ _03925_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06218_ _01129_ _01094_ _01134_ _01141_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__a211o_1
XFILLER_0_130_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07198_ _01865_ rvsingle.dp.rf.rf\[19\]\[17\] _01626_ _02118_ VGND VGND VPWR VPWR
+ _02119_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06149_ _01067_ _01069_ _01072_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09908_ _04364_ _04141_ _04733_ DataAdr[1] VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__o31a_1
X_09839_ _04398_ _04665_ _04670_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[27\] sky130_fd_sc_hd__o21ai_1
X_12850_ clknet_leaf_40_clk _00308_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _04918_ _04928_ _05417_ _04915_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__nor4b_4
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ clknet_leaf_45_clk _00239_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _05716_ net287 _05817_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__mux2_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11663_ _05788_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13402_ clknet_leaf_5_clk _00830_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10614_ _04790_ net745 _05205_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_927 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11594_ _05757_ net486 _05729_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13333_ clknet_leaf_76_clk rvsingle.dp.PCNext\[10\] _00010_ VGND VGND VPWR VPWR PC[10]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10545_ _05149_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_130_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_130_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13264_ clknet_leaf_67_clk _00722_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10476_ _04828_ net539 _05110_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__mux2_1
X_12215_ _06068_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13195_ clknet_leaf_92_clk _00653_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_12146_ _05769_ _05770_ _06007_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12077_ _06005_ _05973_ _06006_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__o21ai_1
X_11028_ _05354_ net772 _05443_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12979_ clknet_leaf_34_clk _00437_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_16 DataAdr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 Instr[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_38 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _02379_ rvsingle.dp.rf.rf\[7\]\[11\] _02031_ _03090_ VGND VGND VPWR VPWR
+ _03091_ sky130_fd_sc_hd__o211ai_1
XANTENNA_49 ReadData[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07121_ _01383_ rvsingle.dp.rf.rf\[6\]\[18\] VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_121_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07052_ _01634_ _01967_ _01972_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07954_ _02873_ _01848_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__a21oi_1
X_06905_ rvsingle.dp.rf.rf\[24\]\[23\] rvsingle.dp.rf.rf\[25\]\[23\] _01335_ VGND
+ VGND VPWR VPWR _01826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07885_ _01828_ rvsingle.dp.rf.rf\[14\]\[2\] _01299_ VGND VGND VPWR VPWR _02806_
+ sky130_fd_sc_hd__o21a_1
X_09624_ _04472_ _04473_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__xor2_1
X_06836_ _01749_ _01756_ _01526_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09555_ _04397_ _02801_ _04410_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06767_ _01687_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08506_ _03424_ _01111_ _03426_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09486_ _04377_ _01536_ _01577_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__and3_2
XFILLER_0_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06698_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08437_ _01499_ rvsingle.dp.rf.rf\[20\]\[9\] VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08368_ _01694_ _03288_ _01699_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07319_ _01595_ rvsingle.dp.rf.rf\[2\]\[16\] VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_112_clk sky130_fd_sc_hd__clkbuf_16
X_08299_ _03171_ _03218_ _01591_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_144_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10330_ _04834_ rvsingle.dp.rf.rf\[26\]\[19\] _05033_ VGND VGND VPWR VPWR _05042_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10261_ _04834_ _04970_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__nand2_1
X_12000_ _04876_ net262 _05960_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__mux2_1
X_10192_ _04959_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12902_ clknet_leaf_114_clk _00360_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_12833_ clknet_leaf_137_clk _00291_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ clknet_leaf_149_clk _00222_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _05794_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__clkbuf_8
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ clknet_leaf_18_clk _00153_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11646_ _05782_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_103_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_103_clk sky130_fd_sc_hd__clkbuf_16
X_11577_ _04814_ _04973_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13316_ clknet_leaf_131_clk _00774_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10528_ _05158_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold809 rvsingle.dp.rf.rf\[28\]\[7\] VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13247_ clknet_leaf_145_clk _00705_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10459_ net8 _05103_ _05116_ _04970_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13178_ clknet_leaf_20_clk _00636_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12129_ _05757_ net608 _06031_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07670_ rvsingle.dp.rf.rf\[12\]\[5\] rvsingle.dp.rf.rf\[13\]\[5\] rvsingle.dp.rf.rf\[14\]\[5\]
+ rvsingle.dp.rf.rf\[15\]\[5\] _01462_ _01727_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__mux4_1
X_06621_ _01091_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__buf_6
X_09340_ _04252_ _04253_ _04137_ _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__a31oi_4
X_06552_ _01192_ rvsingle.dp.rf.rf\[14\]\[21\] VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09271_ _01181_ _01185_ _01249_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__a21oi_1
X_06483_ _01378_ _01387_ _01391_ _01404_ _01154_ VGND VGND VPWR VPWR WriteData[28]
+ sky130_fd_sc_hd__o311a_4
XFILLER_0_28_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08222_ _03111_ _01870_ _01485_ _03142_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08153_ _03070_ _03071_ _02323_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_126_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07104_ rvsingle.dp.rf.rf\[29\]\[18\] _01861_ _01759_ _02024_ VGND VGND VPWR VPWR
+ _02025_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_70_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08084_ rvsingle.dp.rf.rf\[7\]\[1\] _01606_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07035_ _01461_ _01952_ _01955_ _01447_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08986_ _01189_ _03899_ _03905_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__or3_2
X_07937_ _02847_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07868_ _01148_ rvsingle.dp.rf.rf\[18\]\[2\] _01611_ _02788_ VGND VGND VPWR VPWR
+ _02789_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_98_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06819_ _01581_ _01684_ _01486_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09607_ _04427_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__buf_2
X_07799_ _02364_ _02714_ _02719_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__nand3_1
XFILLER_0_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09538_ _04288_ _04286_ VGND VGND VPWR VPWR DataAdr[28] sky130_fd_sc_hd__nand2_8
XFILLER_0_167_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09469_ PC[0] VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11500_ _05476_ net282 _05695_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12480_ clknet_leaf_118_clk _00964_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11431_ _05664_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11362_ _05626_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13101_ clknet_leaf_44_clk _00559_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ _05021_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__buf_6
XFILLER_0_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11293_ _05295_ net729 _05580_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__mux2_1
X_13032_ clknet_leaf_102_clk _00490_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10244_ _04796_ rvsingle.dp.rf.rf\[27\]\[12\] _04989_ VGND VGND VPWR VPWR _04995_
+ sky130_fd_sc_hd__mux2_1
X_10175_ _04950_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12816_ clknet_leaf_71_clk _00274_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12747_ clknet_leaf_88_clk _00205_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12678_ clknet_leaf_113_clk _00136_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11629_ net140 _05779_ _05735_ _05501_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold606 rvsingle.dp.rf.rf\[17\]\[27\] VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold617 rvsingle.dp.rf.rf\[11\]\[26\] VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold628 rvsingle.dp.rf.rf\[12\]\[18\] VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 rvsingle.dp.rf.rf\[27\]\[2\] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _02150_ _01482_ _01486_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__a21o_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ rvsingle.dp.rf.rf\[7\]\[15\] _02627_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__or2b_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07722_ _02337_ _02639_ _02640_ _01564_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_109_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07653_ _02550_ _02569_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06604_ rvsingle.dp.rf.rf\[23\]\[21\] _01509_ _01524_ VGND VGND VPWR VPWR _01525_
+ sky130_fd_sc_hd__o21ai_1
X_07584_ _01152_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09323_ _03830_ _04238_ _03827_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06535_ _01455_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09254_ _04171_ _03772_ _01927_ _04172_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06466_ rvsingle.dp.rf.rf\[16\]\[28\] rvsingle.dp.rf.rf\[17\]\[28\] rvsingle.dp.rf.rf\[18\]\[28\]
+ rvsingle.dp.rf.rf\[19\]\[28\] _01139_ _01107_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08205_ _01295_ rvsingle.dp.rf.rf\[23\]\[11\] _01808_ _03125_ VGND VGND VPWR VPWR
+ _03126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09185_ _01128_ rvsingle.dp.rf.rf\[0\]\[31\] VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06397_ _01195_ rvsingle.dp.rf.rf\[12\]\[29\] VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08136_ _02469_ _02608_ _02666_ _02664_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08067_ _01207_ _02987_ _02447_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_102_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07018_ rvsingle.dp.rf.rf\[28\]\[19\] rvsingle.dp.rf.rf\[29\]\[19\] _01691_ VGND
+ VGND VPWR VPWR _01939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08969_ rvsingle.dp.rf.rf\[24\]\[25\] rvsingle.dp.rf.rf\[25\]\[25\] rvsingle.dp.rf.rf\[26\]\[25\]
+ rvsingle.dp.rf.rf\[27\]\[25\] _01330_ _01302_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__mux4_1
X_11980_ _05344_ net386 _05949_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10931_ _05391_ rvsingle.dp.rf.rf\[18\]\[14\] _05387_ VGND VGND VPWR VPWR _05392_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10862_ _05337_ _05338_ _05339_ _05084_ net205 VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__o41a_1
XFILLER_0_79_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12601_ clknet_leaf_7_clk _00059_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ _04877_ net591 _05298_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12532_ clknet_leaf_62_clk _01016_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12463_ clknet_leaf_39_clk _00947_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11414_ _05655_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__clkbuf_1
X_12394_ clknet_leaf_83_clk _00878_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11345_ _05617_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11276_ _05568_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__buf_6
X_13015_ clknet_leaf_11_clk _00473_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10227_ _04760_ rvsingle.dp.rf.rf\[27\]\[4\] _04978_ VGND VGND VPWR VPWR _04986_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10158_ _04790_ net434 _04941_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 rvsingle.dp.rf.rf\[1\]\[9\] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlygate4sd3_1
X_10089_ _04879_ _04880_ _04881_ ReadData[28] _04715_ VGND VGND VPWR VPWR _04888_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_18_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06320_ _01197_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06251_ Instr[6] Instr[3] Instr[2] VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__nand3_2
XFILLER_0_115_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06182_ _01105_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold403 rvsingle.dp.rf.rf\[2\]\[16\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold414 rvsingle.dp.rf.rf\[6\]\[18\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold425 rvsingle.dp.rf.rf\[26\]\[25\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold436 rvsingle.dp.rf.rf\[24\]\[21\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold447 rvsingle.dp.rf.rf\[20\]\[30\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 rvsingle.dp.rf.rf\[14\]\[25\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 rvsingle.dp.rf.rf\[26\]\[8\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _04364_ _04430_ _04431_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _04398_ _04692_ _04700_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[30\] sky130_fd_sc_hd__o21ai_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _03742_ _03743_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nor2_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _01513_ rvsingle.dp.rf.rf\[10\]\[15\] _02059_ _03674_ VGND VGND VPWR VPWR
+ _03675_ sky130_fd_sc_hd__o211a_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _01797_ rvsingle.dp.rf.rf\[0\]\[5\] VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08685_ rvsingle.dp.rf.rf\[27\]\[14\] _01487_ _03605_ VGND VGND VPWR VPWR _03606_
+ sky130_fd_sc_hd__o21ai_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_92_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ rvsingle.dp.rf.rf\[25\]\[4\] _01295_ _01308_ _02556_ VGND VGND VPWR VPWR
+ _02557_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_166_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07567_ _01110_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__buf_8
XFILLER_0_165_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09306_ _04221_ _04159_ _04161_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__o21bai_4
X_06518_ rvsingle.dp.rf.rf\[21\]\[21\] _01296_ _01437_ _01438_ VGND VGND VPWR VPWR
+ _01439_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07498_ _01552_ _02415_ _02416_ _02329_ _02418_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_63_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09237_ _04154_ _04155_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__nor2_2
XFILLER_0_35_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06449_ rvsingle.dp.rf.rf\[14\]\[28\] rvsingle.dp.rf.rf\[15\]\[28\] _01194_ VGND
+ VGND VPWR VPWR _01371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09168_ rvsingle.dp.rf.rf\[24\]\[31\] rvsingle.dp.rf.rf\[25\]\[31\] rvsingle.dp.rf.rf\[26\]\[31\]
+ rvsingle.dp.rf.rf\[27\]\[31\] _02212_ _01120_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08119_ _03036_ _03037_ _01502_ _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_43_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09099_ _01138_ rvsingle.dp.rf.rf\[6\]\[26\] _03840_ VGND VGND VPWR VPWR _04019_
+ sky130_fd_sc_hd__o21ai_1
X_11130_ _05500_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11061_ _05113_ _05114_ _05115_ _05061_ _04769_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10012_ _04564_ _04565_ _04364_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11963_ _05740_ net314 _05940_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10914_ _05381_ net491 _05373_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11894_ _05910_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10845_ _05337_ _05338_ _05339_ _05084_ net184 VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__o41a_1
XFILLER_0_27_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10776_ _05295_ net685 _05285_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12515_ clknet_leaf_127_clk _00999_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12446_ clknet_leaf_135_clk _00930_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12377_ clknet_leaf_17_clk _00861_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11328_ _05322_ net473 _05607_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11259_ _05571_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
X_08470_ rvsingle.dp.rf.rf\[19\]\[9\] _02303_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07421_ rvsingle.dp.rf.rf\[7\]\[7\] _01557_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__or2b_1
XFILLER_0_148_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07352_ _01172_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__buf_6
XFILLER_0_128_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06303_ _01203_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__buf_4
XFILLER_0_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07283_ _01722_ _02201_ _02203_ _01478_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_61_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09022_ _01089_ rvsingle.dp.rf.rf\[19\]\[27\] _03941_ VGND VGND VPWR VPWR _03942_
+ sky130_fd_sc_hd__o21a_1
X_06234_ rvsingle.dp.rf.rf\[16\]\[30\] rvsingle.dp.rf.rf\[17\]\[30\] rvsingle.dp.rf.rf\[18\]\[30\]
+ rvsingle.dp.rf.rf\[19\]\[30\] _01128_ _01107_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold200 rvsingle.dp.rf.rf\[19\]\[22\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
X_06165_ _01088_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold211 rvsingle.dp.rf.rf\[3\]\[6\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 rvsingle.dp.rf.rf\[12\]\[29\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold233 rvsingle.dp.rf.rf\[2\]\[30\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 rvsingle.dp.rf.rf\[1\]\[24\] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 rvsingle.dp.rf.rf\[11\]\[29\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold266 rvsingle.dp.rf.rf\[23\]\[30\] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 rvsingle.dp.rf.rf\[7\]\[28\] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 rvsingle.dp.rf.rf\[8\]\[29\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09924_ _04748_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__clkbuf_1
Xhold299 rvsingle.dp.rf.rf\[11\]\[27\] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _04618_ PC[28] _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__a21o_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08806_ _01338_ _01201_ _01245_ _03713_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__o311a_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06998_ _01915_ _01916_ _01918_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__o21ai_1
X_09786_ _04618_ PC[22] _04619_ _04620_ _04621_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__a221o_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ rvsingle.dp.rf.rf\[21\]\[15\] _01877_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__or2b_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_106 _01247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_117 _01433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _01499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ rvsingle.dp.rf.rf\[16\]\[14\] rvsingle.dp.rf.rf\[17\]\[14\] rvsingle.dp.rf.rf\[18\]\[14\]
+ rvsingle.dp.rf.rf\[19\]\[14\] _01426_ _02162_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__mux4_1
XANTENNA_139 _01558_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _02537_ _02539_ _02273_ _01217_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__a31oi_2
X_08599_ rvsingle.dp.rf.rf\[13\]\[12\] _01618_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__and2b_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10630_ _05215_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10561_ _04840_ net669 _05151_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12300_ _04746_ rvsingle.dp.rf.rf\[30\]\[2\] _06099_ VGND VGND VPWR VPWR _06101_
+ sky130_fd_sc_hd__mux2_1
X_13280_ clknet_leaf_13_clk _00738_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10492_ _04870_ net678 _05126_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12231_ _06069_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12162_ _05004_ _05328_ _06052_ net211 VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11113_ _05318_ net795 _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12093_ _04769_ rvsingle.dp.rf.rf\[0\]\[6\] _06010_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__mux2_1
X_11044_ _05454_ _05415_ _05455_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12995_ clknet_leaf_116_clk _00453_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11946_ _05721_ _05937_ _05938_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _04738_ _04733_ _05835_ _04739_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__or4b_2
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10828_ _05085_ _05328_ _05325_ net210 VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10759_ _05286_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12429_ clknet_leaf_45_clk _00913_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07970_ rvsingle.dp.rf.rf\[24\]\[0\] _02005_ _01530_ VGND VGND VPWR VPWR _02891_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06921_ _01645_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06852_ _01761_ _01765_ _01634_ _01772_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__o211ai_2
X_09640_ _04484_ _04486_ _04488_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09571_ _04425_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__buf_6
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06783_ rvsingle.dp.rf.rf\[0\]\[20\] rvsingle.dp.rf.rf\[1\]\[20\] rvsingle.dp.rf.rf\[2\]\[20\]
+ rvsingle.dp.rf.rf\[3\]\[20\] _01469_ _01471_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_47_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
X_08522_ rvsingle.dp.rf.rf\[3\]\[13\] _01752_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08453_ _01711_ _03368_ _03373_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07404_ _01630_ rvsingle.dp.rf.rf\[14\]\[7\] _01259_ _02324_ VGND VGND VPWR VPWR
+ _02325_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_92_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08384_ rvsingle.dp.rf.rf\[20\]\[8\] rvsingle.dp.rf.rf\[21\]\[8\] _01191_ VGND VGND
+ VPWR VPWR _03305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07335_ _02239_ _02244_ _01378_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_61_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07266_ rvsingle.dp.rf.rf\[16\]\[16\] rvsingle.dp.rf.rf\[17\]\[16\] _01417_ VGND
+ VGND VPWR VPWR _02187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09005_ _01193_ rvsingle.dp.rf.rf\[8\]\[27\] VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06217_ _01090_ rvsingle.dp.rf.rf\[15\]\[30\] _01107_ _01140_ VGND VGND VPWR VPWR
+ _01141_ sky130_fd_sc_hd__o211a_1
X_07197_ _02117_ rvsingle.dp.rf.rf\[18\]\[17\] VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06148_ _01071_ _01061_ _01062_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09907_ _04732_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__clkbuf_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _04366_ _04668_ _04669_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__nand3_1
XFILLER_0_38_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09769_ _04589_ _04604_ _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__a21oi_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _05858_ _05831_ _05859_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__o21ai_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ clknet_leaf_51_clk _00238_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11731_ _05825_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__clkbuf_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11662_ _05716_ net285 _05775_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13401_ clknet_leaf_32_clk _00829_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10613_ _05193_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__buf_8
X_11593_ _04858_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10544_ _05166_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__clkbuf_1
X_13332_ clknet_leaf_74_clk rvsingle.dp.PCNext\[9\] _00009_ VGND VGND VPWR VPWR PC[9]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13263_ clknet_leaf_48_clk _00721_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10475_ _05124_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12214_ _06068_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__inv_2
X_13194_ clknet_leaf_102_clk _00652_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_12145_ net61 VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12076_ _05769_ _05770_ _05973_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__o21ai_1
X_11027_ _05446_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12978_ clknet_leaf_40_clk _00436_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11929_ _04869_ net260 _05924_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_17 DataAdr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_28 Instr[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 ReadData[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07120_ _02027_ _02040_ _01682_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__nand3_4
XFILLER_0_55_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07051_ _01969_ _01632_ _01971_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07953_ rvsingle.dp.rf.rf\[10\]\[0\] _01493_ _01552_ VGND VGND VPWR VPWR _02874_
+ sky130_fd_sc_hd__o21ai_1
X_06904_ rvsingle.dp.rf.rf\[28\]\[23\] rvsingle.dp.rf.rf\[29\]\[23\] rvsingle.dp.rf.rf\[30\]\[23\]
+ rvsingle.dp.rf.rf\[31\]\[23\] _01463_ _01471_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07884_ rvsingle.dp.rf.rf\[13\]\[2\] _01440_ _02268_ _02804_ VGND VGND VPWR VPWR
+ _02805_ sky130_fd_sc_hd__o211ai_1
X_09623_ Instr[28] PC[8] _04465_ _04466_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__o2bb2a_1
X_06835_ _01565_ _01751_ _01755_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__nand3_1
X_09554_ _04397_ _02801_ _04371_ _04399_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__a2bb2oi_2
X_06766_ _01293_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__buf_4
XFILLER_0_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08505_ rvsingle.dp.rf.rf\[23\]\[13\] _01860_ _03425_ VGND VGND VPWR VPWR _03426_
+ sky130_fd_sc_hd__o21ai_1
X_09485_ _04383_ VGND VGND VPWR VPWR WriteData[22] sky130_fd_sc_hd__clkbuf_4
X_06697_ _01135_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08436_ _01619_ rvsingle.dp.rf.rf\[18\]\[9\] _01620_ _03356_ VGND VGND VPWR VPWR
+ _03357_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08367_ rvsingle.dp.rf.rf\[0\]\[8\] rvsingle.dp.rf.rf\[1\]\[8\] rvsingle.dp.rf.rf\[2\]\[8\]
+ rvsingle.dp.rf.rf\[3\]\[8\] _01730_ _01808_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__mux4_1
X_07318_ _02235_ _01093_ _02236_ _02238_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08298_ _02473_ _02318_ _03171_ _03218_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07249_ _01420_ rvsingle.dp.rf.rf\[30\]\[17\] VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10260_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_942 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10191_ _04886_ net394 _04952_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12901_ clknet_leaf_108_clk _00359_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ clknet_leaf_115_clk _00290_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12763_ clknet_leaf_142_clk _00221_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _05816_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__clkbuf_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ clknet_leaf_26_clk _00152_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11645_ _05439_ rvsingle.dp.rf.rf\[19\]\[18\] _05775_ VGND VGND VPWR VPWR _05782_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11576_ _05167_ _05748_ _05731_ net172 VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13315_ clknet_leaf_126_clk _00773_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10527_ _04760_ net671 _05152_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13246_ clknet_leaf_147_clk _00704_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10458_ _05113_ _05114_ _05115_ _04924_ _04781_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__o311a_1
XFILLER_0_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13177_ clknet_leaf_16_clk _00635_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10389_ _05076_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__clkbuf_1
X_12128_ _06034_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12059_ _05997_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__clkbuf_1
X_06620_ rvsingle.dp.rf.rf\[15\]\[21\] _01540_ _01260_ VGND VGND VPWR VPWR _01541_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_931 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06551_ rvsingle.dp.rf.rf\[8\]\[21\] rvsingle.dp.rf.rf\[9\]\[21\] rvsingle.dp.rf.rf\[10\]\[21\]
+ rvsingle.dp.rf.rf\[11\]\[21\] _01469_ _01471_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09270_ _04063_ _04137_ _04186_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__nand3_2
XFILLER_0_118_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06482_ _01118_ _01397_ _01403_ _01378_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08221_ _01483_ _02260_ _01177_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__o21a_4
XFILLER_0_117_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08152_ rvsingle.dp.rf.rf\[23\]\[11\] _01539_ _03072_ VGND VGND VPWR VPWR _03073_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07103_ _01097_ rvsingle.dp.rf.rf\[28\]\[18\] VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08083_ _01642_ rvsingle.dp.rf.rf\[4\]\[1\] _03003_ _01667_ VGND VGND VPWR VPWR _03004_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_15_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_944 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07034_ rvsingle.dp.rf.rf\[3\]\[19\] _01441_ _01954_ VGND VGND VPWR VPWR _01955_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ _02191_ _03900_ _03904_ _01219_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07936_ _02803_ _02851_ _02856_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_74_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07867_ rvsingle.dp.rf.rf\[19\]\[2\] _01096_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__or2b_1
XFILLER_0_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09606_ _04456_ _04457_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06818_ _01685_ _01737_ _01738_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07798_ _02031_ _02715_ _02716_ _01502_ _02718_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__o311ai_1
X_09537_ _04199_ _04201_ VGND VGND VPWR VPWR DataAdr[27] sky130_fd_sc_hd__nand2_8
XFILLER_0_167_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06749_ _01665_ _01666_ _01668_ _01669_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09468_ _01058_ _04367_ _04374_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08419_ _01634_ _03334_ _03339_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__nand3_1
XFILLER_0_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09399_ _02317_ _02377_ _02373_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11430_ _05476_ net611 _05657_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11361_ _05439_ net618 _05618_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13100_ clknet_leaf_53_clk _00558_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10312_ _05032_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__clkbuf_1
X_11292_ _05588_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13031_ clknet_leaf_101_clk _00489_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10243_ _04994_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_783 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10174_ _04834_ net732 _04941_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12815_ clknet_leaf_27_clk _00273_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ clknet_leaf_81_clk _00204_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12677_ clknet_leaf_114_clk _00135_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11628_ net204 _05779_ _05734_ _05501_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11559_ _04773_ _05732_ _05733_ _05097_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__and4_1
Xhold607 rvsingle.dp.rf.rf\[8\]\[2\] VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold618 rvsingle.dp.rf.rf\[14\]\[18\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold629 rvsingle.dp.rf.rf\[0\]\[4\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13229_ clknet_leaf_90_clk _00687_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ rvsingle.dp.rf.rf\[5\]\[15\] _01602_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__and2b_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07721_ _01797_ rvsingle.dp.rf.rf\[26\]\[5\] _01647_ _02641_ VGND VGND VPWR VPWR
+ _02642_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07652_ _02570_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__nand2_1
X_06603_ _01493_ rvsingle.dp.rf.rf\[22\]\[21\] _01523_ VGND VGND VPWR VPWR _01524_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07583_ _02484_ _02492_ _01377_ _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_149_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09322_ _04165_ _04237_ _03774_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__a21oi_1
X_06534_ _01454_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__buf_8
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09253_ _04168_ _04169_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__nand2_1
X_06465_ _01113_ _01379_ _01386_ _01118_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08204_ _01725_ rvsingle.dp.rf.rf\[22\]\[11\] VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09184_ rvsingle.dp.rf.rf\[2\]\[31\] rvsingle.dp.rf.rf\[3\]\[31\] _01100_ VGND VGND
+ VPWR VPWR _04104_ sky130_fd_sc_hd__mux2_1
X_06396_ rvsingle.dp.rf.rf\[8\]\[29\] rvsingle.dp.rf.rf\[9\]\[29\] rvsingle.dp.rf.rf\[10\]\[29\]
+ rvsingle.dp.rf.rf\[11\]\[29\] _01195_ _01202_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08135_ _03055_ _02572_ _02570_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__nand3_2
XFILLER_0_70_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08066_ rvsingle.dp.rf.rf\[20\]\[1\] rvsingle.dp.rf.rf\[21\]\[1\] rvsingle.dp.rf.rf\[22\]\[1\]
+ rvsingle.dp.rf.rf\[23\]\[1\] _02440_ _01470_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07017_ _01441_ rvsingle.dp.rf.rf\[31\]\[19\] _01301_ _01937_ VGND VGND VPWR VPWR
+ _01938_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08968_ rvsingle.dp.rf.rf\[28\]\[25\] rvsingle.dp.rf.rf\[29\]\[25\] rvsingle.dp.rf.rf\[30\]\[25\]
+ rvsingle.dp.rf.rf\[31\]\[25\] _01194_ _01303_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__mux4_1
X_07919_ _02275_ rvsingle.dp.rf.rf\[27\]\[2\] _02162_ _02839_ VGND VGND VPWR VPWR
+ _02840_ sky130_fd_sc_hd__o211a_1
X_08899_ _01828_ rvsingle.dp.rf.rf\[14\]\[24\] VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__or2_1
X_10930_ _04807_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10861_ _05085_ _05348_ _05325_ net169 VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_168_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12600_ clknet_leaf_33_clk _00058_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10792_ _05305_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12531_ clknet_leaf_32_clk _01015_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12462_ clknet_leaf_72_clk _00946_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11413_ _05428_ net484 _05646_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12393_ clknet_leaf_92_clk _00877_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11344_ _05385_ rvsingle.dp.rf.rf\[14\]\[10\] _05607_ VGND VGND VPWR VPWR _05617_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11275_ _05579_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13014_ clknet_leaf_25_clk _00472_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10226_ net42 _04978_ _04984_ _04985_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__a22o_1
X_10157_ _04929_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__buf_6
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 rvsingle.dp.rf.rf\[1\]\[0\] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10088_ _04887_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12729_ clknet_leaf_8_clk _00187_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06250_ Instr[1] Instr[0] VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06181_ _01104_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold404 rvsingle.dp.rf.rf\[29\]\[9\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold415 rvsingle.dp.rf.rf\[28\]\[14\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 rvsingle.dp.rf.rf\[31\]\[30\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 rvsingle.dp.rf.rf\[2\]\[20\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 rvsingle.dp.rf.rf\[17\]\[9\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 rvsingle.dp.rf.rf\[14\]\[29\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09940_ DataAdr[5] ReadData[5] _04751_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _04366_ _04698_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__nand3_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _03728_ _03699_ _03727_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ rvsingle.dp.rf.rf\[11\]\[15\] _01136_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07704_ _02623_ _02624_ _01111_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__o21ai_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _01613_ rvsingle.dp.rf.rf\[26\]\[14\] _01551_ VGND VGND VPWR VPWR _03605_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ _01191_ rvsingle.dp.rf.rf\[24\]\[4\] VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07566_ rvsingle.dp.rf.rf\[5\]\[4\] _01677_ _02485_ _02486_ VGND VGND VPWR VPWR _02487_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_49_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09305_ _03231_ _03406_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__or2_1
X_06517_ _01192_ rvsingle.dp.rf.rf\[20\]\[21\] VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07497_ _01658_ rvsingle.dp.rf.rf\[2\]\[6\] _01654_ _02417_ VGND VGND VPWR VPWR _02418_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_119_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09236_ _03056_ _02576_ _02661_ _02667_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__nand4_1
X_06448_ rvsingle.dp.rf.rf\[13\]\[28\] _01298_ _01311_ _01369_ VGND VGND VPWR VPWR
+ _01370_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06379_ _01300_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__buf_4
X_09167_ _01219_ _04079_ _01317_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08118_ _02005_ rvsingle.dp.rf.rf\[30\]\[1\] _01104_ _03038_ VGND VGND VPWR VPWR
+ _03039_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09098_ rvsingle.dp.rf.rf\[7\]\[26\] VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__inv_2
X_08049_ _01690_ rvsingle.dp.rf.rf\[8\]\[1\] VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__or2_1
X_11060_ _05463_ net159 _05159_ _05464_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__a22o_1
X_10011_ _04751_ _04256_ _04820_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11962_ _05947_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10913_ _04773_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__buf_2
X_11893_ _05740_ net433 _05902_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10844_ _04965_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10775_ _04833_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__buf_2
X_12514_ clknet_leaf_128_clk _00998_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12445_ clknet_leaf_143_clk _00929_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12376_ clknet_leaf_18_clk _00860_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11327_ _05608_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11258_ _05322_ rvsingle.dp.rf.rf\[15\]\[2\] _05569_ VGND VGND VPWR VPWR _05571_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10209_ _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__buf_1
X_11189_ _05532_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07420_ rvsingle.dp.rf.rf\[5\]\[7\] _01136_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07351_ rvsingle.dp.rf.rf\[15\]\[7\] _02271_ _01300_ VGND VGND VPWR VPWR _02272_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06302_ _01195_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__buf_4
X_07282_ rvsingle.dp.rf.rf\[3\]\[16\] _01296_ _02202_ VGND VGND VPWR VPWR _02203_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09021_ _01098_ rvsingle.dp.rf.rf\[18\]\[27\] _01626_ VGND VGND VPWR VPWR _03941_
+ sky130_fd_sc_hd__o21a_1
X_06233_ _01156_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__buf_8
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06164_ _01087_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__clkbuf_8
Xhold201 rvsingle.dp.rf.rf\[3\]\[13\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 rvsingle.dp.rf.rf\[9\]\[27\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 rvsingle.dp.rf.rf\[2\]\[26\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold234 rvsingle.dp.rf.rf\[25\]\[22\] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 rvsingle.dp.rf.rf\[25\]\[23\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 rvsingle.dp.rf.rf\[23\]\[23\] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold267 rvsingle.dp.rf.rf\[0\]\[30\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 rvsingle.dp.rf.rf\[4\]\[21\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _04747_ rvsingle.dp.rf.rf\[2\]\[2\] _04741_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__mux2_1
Xhold289 rvsingle.dp.rf.rf\[27\]\[28\] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _04618_ PC[28] _04674_ _04676_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__o22a_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _01316_ _03719_ _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__nand3_4
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _04609_ _04606_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__nor2_1
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ _01461_ _01917_ _01447_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__o21a_1
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ rvsingle.dp.rf.rf\[23\]\[15\] _02478_ _01490_ VGND VGND VPWR VPWR _03657_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _01247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _01433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _02093_ _03587_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _01687_ rvsingle.dp.rf.rf\[15\]\[4\] _01708_ _02538_ VGND VGND VPWR VPWR
+ _02539_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_166_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _01630_ rvsingle.dp.rf.rf\[12\]\[12\] VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07549_ _01450_ _02449_ _02462_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10560_ _05167_ _05175_ _05155_ net94 VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_118_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09219_ _04133_ _04116_ _04134_ _04137_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__o211ai_4
X_10491_ net23 _05103_ _05133_ _04970_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12230_ _06069_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12161_ net100 _06052_ _05327_ _04985_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11112_ _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__buf_8
X_12092_ _06015_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__clkbuf_1
Xhold790 rvsingle.dp.rf.rf\[20\]\[2\] VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd3_1
X_11043_ _05364_ _05365_ _05415_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_12994_ clknet_leaf_141_clk _00452_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11945_ _05099_ _05832_ net116 VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11876_ _05721_ _05899_ _05900_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__a21oi_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10827_ _04982_ _04983_ _04981_ _04769_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__or4b_1
XFILLER_0_95_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10758_ _04790_ rvsingle.dp.rf.rf\[20\]\[11\] _05285_ VGND VGND VPWR VPWR _05286_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10689_ _05207_ net423 _05246_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12428_ clknet_leaf_50_clk _00912_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12359_ _06131_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06920_ _01666_ rvsingle.dp.rf.rf\[14\]\[22\] VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__nor2_1
X_06851_ _01655_ _01766_ _01767_ _01768_ _01771_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__o311ai_2
X_09570_ _01080_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__buf_4
X_06782_ _01702_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__clkbuf_8
X_08521_ rvsingle.dp.rf.rf\[1\]\[13\] _01498_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08452_ _03370_ _02291_ _03372_ _01217_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_147_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07403_ rvsingle.dp.rf.rf\[15\]\[7\] _01544_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__or2b_1
XFILLER_0_148_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08383_ rvsingle.dp.rf.rf\[16\]\[8\] rvsingle.dp.rf.rf\[17\]\[8\] rvsingle.dp.rf.rf\[18\]\[8\]
+ rvsingle.dp.rf.rf\[19\]\[8\] _01730_ _01808_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07334_ _02236_ _02249_ _02254_ _01506_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_116_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07265_ rvsingle.dp.rf.rf\[19\]\[16\] _01943_ _02185_ VGND VGND VPWR VPWR _02186_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09004_ net212 VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06216_ _01139_ rvsingle.dp.rf.rf\[14\]\[30\] VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__or2_1
X_07196_ _01752_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__buf_6
X_06147_ _01070_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09906_ net825 VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _04651_ _04666_ _04667_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__nand3_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ PC[20] PC[21] _04590_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__o21a_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _01545_ rvsingle.dp.rf.rf\[6\]\[14\] _02337_ _03639_ VGND VGND VPWR VPWR
+ _03640_ sky130_fd_sc_hd__o211ai_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ PC[14] PC[15] _04522_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__and3_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11730_ _05763_ net281 _05817_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__mux2_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11661_ _05787_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__clkbuf_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13400_ clknet_leaf_24_clk _00828_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10612_ _05204_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11592_ net76 _05726_ _05756_ _05737_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13331_ clknet_leaf_74_clk rvsingle.dp.PCNext\[8\] _00008_ VGND VGND VPWR VPWR PC[8]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_146_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10543_ _04796_ net592 _05151_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13262_ clknet_leaf_53_clk _00720_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10474_ _04824_ net738 _05110_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12213_ _06068_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13193_ clknet_leaf_100_clk _00651_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12144_ _06042_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12075_ net49 VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__inv_2
X_11026_ _05352_ rvsingle.dp.rf.rf\[31\]\[23\] _05443_ VGND VGND VPWR VPWR _05446_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ clknet_leaf_40_clk _00435_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11928_ _05928_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11859_ _05891_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 DataAdr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_29 Instr[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07050_ rvsingle.dp.rf.rf\[23\]\[19\] _01842_ _01970_ VGND VGND VPWR VPWR _01971_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07952_ net248 VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__inv_2
X_06903_ _01722_ _01823_ _01218_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__o21ai_1
X_07883_ _01419_ rvsingle.dp.rf.rf\[12\]\[2\] VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__or2_1
X_09622_ _04470_ _04471_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__nor2_1
X_06834_ _01646_ rvsingle.dp.rf.rf\[9\]\[23\] _01754_ VGND VGND VPWR VPWR _01755_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09553_ _04407_ _04408_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__and2b_1
X_06765_ rvsingle.dp.rf.rf\[8\]\[20\] rvsingle.dp.rf.rf\[9\]\[20\] rvsingle.dp.rf.rf\[10\]\[20\]
+ rvsingle.dp.rf.rf\[11\]\[20\] _01463_ _01471_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08504_ _01544_ rvsingle.dp.rf.rf\[22\]\[13\] _01258_ VGND VGND VPWR VPWR _03425_
+ sky130_fd_sc_hd__o21a_1
X_09484_ _01154_ _01869_ _01896_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__and3_2
X_06696_ _01110_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__buf_8
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08435_ rvsingle.dp.rf.rf\[19\]\[9\] _03258_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__or2b_1
XFILLER_0_109_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08366_ _03284_ _01309_ _01422_ _03286_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_117_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07317_ _01269_ rvsingle.dp.rf.rf\[6\]\[16\] _01491_ _02237_ VGND VGND VPWR VPWR
+ _02238_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08297_ _02505_ _03194_ _03217_ _01083_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__nand4_4
XFILLER_0_6_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07248_ rvsingle.dp.rf.rf\[28\]\[17\] rvsingle.dp.rf.rf\[29\]\[17\] _01432_ VGND
+ VGND VPWR VPWR _02169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07179_ _02097_ _02066_ _02068_ _02099_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_30_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10190_ _04958_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__clkbuf_1
X_12900_ clknet_leaf_110_clk _00358_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12831_ clknet_leaf_16_clk _00289_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ clknet_leaf_4_clk _00220_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11713_ _05398_ rvsingle.dp.rf.rf\[10\]\[20\] _05806_ VGND VGND VPWR VPWR _05816_
+ sky130_fd_sc_hd__mux2_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ clknet_leaf_60_clk _00151_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ net199 _05778_ _05751_ _05457_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11575_ _04976_ _05417_ _04807_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__or3b_2
X_13314_ clknet_leaf_120_clk _00772_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10526_ net150 _05155_ _05156_ _05157_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13245_ clknet_leaf_136_clk _00703_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10457_ _04880_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13176_ clknet_leaf_22_clk _00634_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_10388_ _04790_ rvsingle.dp.rf.rf\[25\]\[11\] _05071_ VGND VGND VPWR VPWR _05076_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12127_ _04852_ net398 _06031_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12058_ _04852_ net527 _05994_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__mux2_1
X_11009_ _05436_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_943 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06550_ _01470_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__clkbuf_8
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06481_ _01134_ _01398_ _01400_ _01402_ _01118_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_290 _05004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08220_ _03112_ _03140_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08151_ _01498_ rvsingle.dp.rf.rf\[22\]\[11\] _01519_ VGND VGND VPWR VPWR _03072_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07102_ rvsingle.dp.rf.rf\[31\]\[18\] _01865_ _01655_ VGND VGND VPWR VPWR _02023_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08082_ rvsingle.dp.rf.rf\[5\]\[1\] _01606_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07033_ _01726_ rvsingle.dp.rf.rf\[2\]\[19\] _01953_ VGND VGND VPWR VPWR _01954_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08984_ _03901_ _01310_ _01230_ _03903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__a211o_1
X_07935_ _02853_ _02854_ _02855_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__nand3_4
X_07866_ rvsingle.dp.rf.rf\[17\]\[2\] _01594_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__and2b_1
X_09605_ PC[7] _04444_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__nor2_1
X_06817_ _01587_ _01684_ _01486_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07797_ _01743_ rvsingle.dp.rf.rf\[6\]\[3\] _01647_ _02717_ VGND VGND VPWR VPWR _02718_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09536_ _04234_ VGND VGND VPWR VPWR DataAdr[26] sky130_fd_sc_hd__clkinv_4
X_06748_ _01256_ rvsingle.dp.rf.rf\[22\]\[20\] VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09467_ _04370_ _04373_ _04366_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__o21ai_1
X_06679_ _01599_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08418_ _01105_ _03335_ _03336_ _02488_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09398_ _04311_ _02464_ _04310_ _04125_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__a31o_1
XFILLER_0_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08349_ rvsingle.dp.rf.rf\[17\]\[8\] _03258_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11360_ _05625_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__clkbuf_1
X_10311_ _04786_ net315 _05022_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11291_ _05439_ rvsingle.dp.rf.rf\[15\]\[18\] _05580_ VGND VGND VPWR VPWR _05588_
+ sky130_fd_sc_hd__mux2_1
X_13030_ clknet_leaf_112_clk _00488_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10242_ _04790_ rvsingle.dp.rf.rf\[27\]\[11\] _04989_ VGND VGND VPWR VPWR _04994_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10173_ _04949_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12814_ clknet_leaf_70_clk _00272_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ clknet_leaf_96_clk _00203_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ clknet_leaf_107_clk _00134_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11627_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11558_ net60 _05731_ _05738_ _05737_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__a22o_1
Xhold608 rvsingle.dp.rf.rf\[0\]\[23\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ _04879_ _04881_ _04880_ _05057_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__o31a_4
XFILLER_0_100_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold619 rvsingle.dp.rf.rf\[21\]\[23\] VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ _05696_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13228_ clknet_leaf_93_clk _00686_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ clknet_leaf_99_clk _00617_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ rvsingle.dp.rf.rf\[27\]\[5\] _01606_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__or2b_1
X_07651_ _02473_ _02318_ _01537_ _02571_ _02530_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06602_ _01489_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__buf_6
X_07582_ _01503_ _02497_ _02502_ _01116_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__o211ai_4
X_09321_ _01931_ _02101_ _02184_ _02265_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__and4_1
XFILLER_0_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06533_ _01197_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09252_ _01836_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06464_ _01380_ _01093_ _01133_ _01385_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08203_ _03114_ _03116_ _01315_ _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09183_ rvsingle.dp.rf.rf\[4\]\[31\] rvsingle.dp.rf.rf\[5\]\[31\] rvsingle.dp.rf.rf\[6\]\[31\]
+ rvsingle.dp.rf.rf\[7\]\[31\] _02212_ _01120_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06395_ _01316_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__buf_8
XFILLER_0_160_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08134_ _02530_ _02533_ _01591_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08065_ _02983_ _01437_ _01702_ _02985_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_141_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07016_ _01695_ rvsingle.dp.rf.rf\[30\]\[19\] VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08967_ _03884_ _01311_ _01231_ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a211oi_2
X_07918_ _01191_ rvsingle.dp.rf.rf\[26\]\[2\] VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__or2_1
X_08898_ rvsingle.dp.rf.rf\[12\]\[24\] rvsingle.dp.rf.rf\[13\]\[24\] _01335_ VGND
+ VGND VPWR VPWR _03819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07849_ rvsingle.dp.rf.rf\[7\]\[2\] _01096_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__or2b_1
XFILLER_0_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10860_ _04834_ _05316_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09519_ _03050_ _03047_ _03051_ _04143_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_149_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10791_ _05304_ net589 _05298_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__mux2_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12530_ clknet_leaf_35_clk _01014_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12461_ clknet_leaf_44_clk _00945_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11412_ _05654_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12392_ clknet_leaf_104_clk _00876_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11343_ _05616_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11274_ _05385_ rvsingle.dp.rf.rf\[15\]\[10\] _05569_ VGND VGND VPWR VPWR _05579_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13013_ clknet_leaf_65_clk _00471_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10225_ _04972_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__buf_6
X_10156_ _04940_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 rvsingle.dp.rf.rf\[25\]\[3\] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _04886_ net391 _04847_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10989_ _05425_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12728_ clknet_leaf_32_clk _00186_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12659_ clknet_leaf_35_clk _00117_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06180_ _01103_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold405 rvsingle.dp.rf.rf\[26\]\[26\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 rvsingle.dp.rf.rf\[26\]\[4\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_868 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold427 rvsingle.dp.rf.rf\[14\]\[28\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold438 rvsingle.dp.rf.rf\[15\]\[12\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold449 rvsingle.dp.rf.rf\[15\]\[28\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _04696_ _04697_ _04693_ _04694_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__nand4_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _03741_ _02261_ _03733_ _03731_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__a211oi_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _03661_ _01146_ _03672_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__nand3_4
X_07703_ rvsingle.dp.rf.rf\[5\]\[5\] _01594_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08683_ rvsingle.dp.rf.rf\[25\]\[14\] _01769_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07634_ _02552_ _02554_ _02273_ _01217_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__a31oi_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07565_ _01136_ rvsingle.dp.rf.rf\[4\]\[4\] VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__or2_1
X_09304_ _03648_ _03650_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__nand2_1
X_06516_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__buf_8
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07496_ rvsingle.dp.rf.rf\[3\]\[6\] _01557_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09235_ _02374_ _02377_ _02464_ _02468_ _02475_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__o2111ai_4
X_06447_ _01338_ rvsingle.dp.rf.rf\[12\]\[28\] VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09166_ _01210_ _04081_ _04083_ _01224_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__o311a_1
XFILLER_0_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06378_ _01299_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08117_ rvsingle.dp.rf.rf\[31\]\[1\] _01124_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__or2b_1
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09097_ _04014_ _01093_ _03782_ _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_142_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08048_ _01440_ rvsingle.dp.rf.rf\[11\]\[1\] _02162_ _02968_ VGND VGND VPWR VPWR
+ _02969_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10010_ _04140_ _04141_ _04732_ ReadData[17] VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__or4b_1
X_09999_ _04228_ _04396_ _04751_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__a21oi_1
X_11961_ _04773_ net549 _05940_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__mux2_1
X_10912_ _05380_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__clkbuf_1
X_11892_ _05909_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10843_ _04917_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__buf_4
XFILLER_0_168_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10774_ _05294_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12513_ clknet_leaf_139_clk _00997_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12444_ clknet_leaf_146_clk _00928_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12375_ clknet_leaf_18_clk _00859_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11326_ _05318_ net701 _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11257_ _05570_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10208_ _04713_ _04919_ _04737_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__and3_1
X_11188_ _05531_ net816 _05528_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__mux2_1
X_10139_ _04747_ net393 _04930_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07350_ _01293_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__buf_4
X_06301_ _01223_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07281_ _01417_ rvsingle.dp.rf.rf\[2\]\[16\] _01244_ VGND VGND VPWR VPWR _02202_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_171_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_151_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_151_clk sky130_fd_sc_hd__clkbuf_16
X_09020_ rvsingle.dp.rf.rf\[16\]\[27\] rvsingle.dp.rf.rf\[17\]\[27\] _01269_ VGND
+ VGND VPWR VPWR _03940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06232_ _01155_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__buf_8
XFILLER_0_5_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06163_ _01086_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold202 rvsingle.dp.rf.rf\[19\]\[15\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 rvsingle.dp.rf.rf\[19\]\[25\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 rvsingle.dp.rf.rf\[3\]\[11\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 rvsingle.dp.rf.rf\[23\]\[28\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold246 rvsingle.dp.rf.rf\[23\]\[14\] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold257 rvsingle.dp.rf.rf\[19\]\[28\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 rvsingle.dp.rf.rf\[30\]\[26\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09922_ _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__clkbuf_2
Xhold279 rvsingle.dp.rf.rf\[28\]\[21\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09853_ PC[29] _04681_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__a21o_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _01461_ _03720_ _03724_ _01218_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__o211ai_2
X_09784_ _04590_ PC[23] VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__or2_1
X_06996_ rvsingle.dp.rf.rf\[12\]\[22\] rvsingle.dp.rf.rf\[13\]\[22\] rvsingle.dp.rf.rf\[14\]\[22\]
+ rvsingle.dp.rf.rf\[15\]\[22\] _01335_ _01199_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__mux4_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _01595_ rvsingle.dp.rf.rf\[22\]\[15\] VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__nor2_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _01247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08666_ rvsingle.dp.rf.rf\[20\]\[14\] rvsingle.dp.rf.rf\[21\]\[14\] rvsingle.dp.rf.rf\[22\]\[14\]
+ rvsingle.dp.rf.rf\[23\]\[14\] _01241_ _01953_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__mux4_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _01690_ rvsingle.dp.rf.rf\[14\]\[4\] VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08597_ _01499_ rvsingle.dp.rf.rf\[10\]\[12\] _02059_ _03517_ VGND VGND VPWR VPWR
+ _03518_ sky130_fd_sc_hd__o211a_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07548_ _01452_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__buf_8
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_142_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_142_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07479_ _02395_ _02396_ _02397_ _01111_ _02399_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_146_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09218_ _04136_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__buf_8
XFILLER_0_91_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10490_ _05113_ _05114_ _05115_ _04924_ _05132_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__o311a_1
XFILLER_0_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09149_ _01232_ _04064_ _04066_ _04068_ _01224_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12160_ _05004_ _05326_ _06052_ net203 VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11111_ _04737_ _04919_ _04733_ _05371_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__or4_4
XFILLER_0_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12091_ _04764_ rvsingle.dp.rf.rf\[0\]\[5\] _06010_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__mux2_1
Xhold780 rvsingle.dp.rf.rf\[23\]\[11\] VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 rvsingle.dp.rf.rf\[0\]\[21\] VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11042_ net81 VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12993_ clknet_leaf_140_clk _00451_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11944_ _04721_ _04920_ _05830_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11875_ net111 _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__nor2_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ _05327_ _05069_ _05068_ _05325_ net13 VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__a32o_1
XFILLER_0_156_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10757_ _05273_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__buf_8
XFILLER_0_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_133_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_133_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10688_ _05247_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12427_ clknet_leaf_64_clk _00911_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12358_ _04903_ net258 _06121_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11309_ _05597_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__clkbuf_1
X_12289_ _06093_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06850_ _01656_ rvsingle.dp.rf.rf\[2\]\[23\] _01660_ _01770_ VGND VGND VPWR VPWR
+ _01771_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06781_ _01172_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__buf_8
X_08520_ _01642_ rvsingle.dp.rf.rf\[0\]\[13\] VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08451_ rvsingle.dp.rf.rf\[15\]\[9\] _01827_ _03371_ VGND VGND VPWR VPWR _03372_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07402_ _01110_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__buf_6
XFILLER_0_147_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08382_ _02093_ _03302_ _01221_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07333_ _02250_ _02251_ _01132_ _02253_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_124_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07264_ _01336_ rvsingle.dp.rf.rf\[18\]\[16\] _01301_ VGND VGND VPWR VPWR _02185_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09003_ _01209_ _03918_ _03922_ _01219_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__o211a_1
X_06215_ _01138_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__buf_8
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07195_ _02114_ _02115_ _01565_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06146_ Instr[1] Instr[0] VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire3 _03143_ VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__buf_2
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09905_ _04121_ _04713_ ReadData[1] _04364_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _04651_ _04666_ _04667_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__a21o_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06979_ _01329_ rvsingle.dp.rf.rf\[18\]\[22\] VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__nor2_1
X_09767_ _04593_ _04600_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__nor2_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ rvsingle.dp.rf.rf\[7\]\[14\] _01877_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__or2b_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ PC[14] _04522_ PC[15] VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _02505_ _03452_ _03429_ _02375_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__a31o_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _05763_ net257 _05775_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__mux2_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10611_ _04786_ net694 _05194_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_115_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_115_clk sky130_fd_sc_hd__clkbuf_16
X_11591_ _04852_ _04968_ _04967_ _05097_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13330_ clknet_leaf_73_clk rvsingle.dp.PCNext\[7\] _00007_ VGND VGND VPWR VPWR PC[7]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10542_ _05165_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13261_ clknet_leaf_90_clk _00719_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10473_ _05123_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12212_ _06068_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13192_ clknet_leaf_121_clk _00650_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12143_ _05639_ net267 _06031_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12074_ _06004_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11025_ _05445_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ clknet_leaf_52_clk _00434_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11927_ _05132_ net249 _05924_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__mux2_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _04876_ net691 _05885_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_106_clk sky130_fd_sc_hd__clkbuf_16
X_10809_ _04725_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_19 DataAdr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11789_ _05853_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07951_ _02868_ _02869_ _01617_ _02871_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06902_ rvsingle.dp.rf.rf\[20\]\[23\] rvsingle.dp.rf.rf\[21\]\[23\] rvsingle.dp.rf.rf\[22\]\[23\]
+ rvsingle.dp.rf.rf\[23\]\[23\] _01463_ _01471_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07882_ _02798_ _02802_ _01485_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__a21oi_4
X_06833_ _01753_ rvsingle.dp.rf.rf\[8\]\[23\] _01604_ VGND VGND VPWR VPWR _01754_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09621_ Instr[29] PC[9] VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__nor2_1
X_09552_ PC[3] _02748_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__nand2_1
X_06764_ _01084_ _01483_ _01591_ _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__o211a_2
X_08503_ _02379_ rvsingle.dp.rf.rf\[21\]\[13\] _03423_ VGND VGND VPWR VPWR _03424_
+ sky130_fd_sc_hd__o21ai_1
X_09483_ _04382_ VGND VGND VPWR VPWR WriteData[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06695_ rvsingle.dp.rf.rf\[13\]\[20\] _01148_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08434_ _03353_ _03354_ _02483_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08365_ _01424_ rvsingle.dp.rf.rf\[7\]\[8\] _01244_ _03285_ VGND VGND VPWR VPWR _03286_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07316_ rvsingle.dp.rf.rf\[7\]\[16\] _01518_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08296_ _03205_ _01682_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__nand3_4
XFILLER_0_117_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07247_ _01478_ _02155_ _02159_ _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07178_ _01223_ _02074_ _02080_ _01317_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09819_ _04590_ PC[26] VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__or2_1
X_12830_ clknet_leaf_0_clk _00288_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ clknet_leaf_32_clk _00219_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _05815_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__clkbuf_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ clknet_leaf_62_clk _00150_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _05471_ _05781_ _05779_ net217 VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11574_ _05167_ _05747_ _05731_ net157 VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_24_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10525_ _05146_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__clkbuf_8
X_13313_ clknet_leaf_132_clk _00771_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13244_ clknet_leaf_12_clk _00702_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10456_ _04881_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13175_ clknet_leaf_65_clk _00633_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10387_ _05075_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__clkbuf_1
X_12126_ _06033_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12057_ _05996_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11008_ _05212_ net812 _05431_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ clknet_leaf_2_clk _00417_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06480_ _01401_ _01093_ _01113_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 _02288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_291 _05004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08150_ rvsingle.dp.rf.rf\[21\]\[11\] _01860_ _01530_ VGND VGND VPWR VPWR _03071_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07101_ _01559_ rvsingle.dp.rf.rf\[30\]\[18\] VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__nor2_1
X_08081_ _02998_ _02999_ _03001_ _01564_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07032_ _01198_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08983_ _01296_ rvsingle.dp.rf.rf\[3\]\[25\] _01434_ _03902_ VGND VGND VPWR VPWR
+ _03903_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07934_ _02473_ _02318_ _01537_ _02698_ _02746_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_138_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07865_ _01847_ rvsingle.dp.rf.rf\[16\]\[2\] VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ PC[5] PC[6] PC[7] _04421_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__and4_2
X_06816_ _01450_ _01714_ _01736_ _01247_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__o211a_4
X_07796_ rvsingle.dp.rf.rf\[7\]\[3\] _01606_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06747_ _01667_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__buf_4
X_09535_ _04249_ VGND VGND VPWR VPWR DataAdr[25] sky130_fd_sc_hd__inv_6
XFILLER_0_149_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09466_ _04371_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06678_ _01130_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08417_ _01513_ rvsingle.dp.rf.rf\[6\]\[9\] _01490_ _03337_ VGND VGND VPWR VPWR _03338_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_136_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09397_ _02464_ _04310_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08348_ _01763_ rvsingle.dp.rf.rf\[16\]\[8\] VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08279_ _01268_ rvsingle.dp.rf.rf\[22\]\[10\] VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10310_ _05031_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11290_ _05587_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10241_ _04993_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__clkbuf_1
X_10172_ _04828_ net707 _04941_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12813_ clknet_leaf_45_clk _00271_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ clknet_leaf_104_clk _00202_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ clknet_leaf_115_clk _00133_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11626_ _05774_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__buf_6
XFILLER_0_108_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11557_ _04769_ _05732_ _05733_ _05097_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold609 rvsingle.dp.rf.rf\[22\]\[20\] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ _05097_ _05058_ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__and3_2
X_11488_ _05334_ net566 _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10439_ _05104_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__clkbuf_1
X_13227_ clknet_leaf_94_clk _00685_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ clknet_leaf_113_clk _00616_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _06024_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__clkbuf_1
X_13089_ clknet_leaf_137_clk _00547_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07650_ Instr[11] _01078_ _02531_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__o21ai_2
X_06601_ _01509_ rvsingle.dp.rf.rf\[21\]\[21\] _01521_ VGND VGND VPWR VPWR _01522_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07581_ _02498_ _02499_ _02500_ _02501_ _02488_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__o221ai_4
X_09320_ _04207_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06532_ _01431_ _01449_ _01450_ _01452_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__a31o_2
XFILLER_0_164_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09251_ _04168_ _04169_ _01927_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__a21boi_1
X_06463_ _01089_ rvsingle.dp.rf.rf\[31\]\[28\] _01106_ _01384_ VGND VGND VPWR VPWR
+ _01385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08202_ _01422_ _03117_ _03122_ _01221_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__o211ai_4
X_09182_ _04100_ _04101_ _01134_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06394_ _01315_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__buf_8
X_08133_ _02751_ _02857_ _02862_ _03053_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_160_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08064_ _02275_ rvsingle.dp.rf.rf\[19\]\[1\] _02162_ _02984_ VGND VGND VPWR VPWR
+ _02985_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07015_ rvsingle.dp.rf.rf\[24\]\[19\] rvsingle.dp.rf.rf\[25\]\[19\] rvsingle.dp.rf.rf\[26\]\[19\]
+ rvsingle.dp.rf.rf\[27\]\[19\] _01469_ _01728_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__mux4_2
XFILLER_0_141_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08966_ _01298_ rvsingle.dp.rf.rf\[19\]\[25\] _01303_ _03885_ VGND VGND VPWR VPWR
+ _03886_ sky130_fd_sc_hd__o211a_1
X_07917_ _02303_ rvsingle.dp.rf.rf\[25\]\[2\] _02837_ VGND VGND VPWR VPWR _02838_
+ sky130_fd_sc_hd__o21a_1
X_08897_ rvsingle.dp.rf.rf\[8\]\[24\] rvsingle.dp.rf.rf\[9\]\[24\] rvsingle.dp.rf.rf\[10\]\[24\]
+ rvsingle.dp.rf.rf\[11\]\[24\] _01463_ _01471_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_95_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
X_07848_ rvsingle.dp.rf.rf\[5\]\[2\] _01492_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__and2b_1
XFILLER_0_151_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07779_ rvsingle.dp.rf.rf\[9\]\[3\] _01087_ _01667_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09518_ _04130_ VGND VGND VPWR VPWR DataAdr[0] sky130_fd_sc_hd__inv_2
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10790_ _04868_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__buf_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09449_ _04153_ _02661_ _04355_ _03058_ _04309_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__a311o_1
XFILLER_0_93_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12460_ clknet_leaf_50_clk _00944_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11411_ _05330_ net726 _05646_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12391_ clknet_leaf_99_clk _00875_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11342_ _05428_ net495 _05607_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11273_ _05578_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13012_ clknet_leaf_61_clk _00470_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10224_ _04981_ _04754_ _04982_ _04983_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__and4b_1
X_10155_ _04786_ rvsingle.dp.rf.rf\[28\]\[10\] _04930_ VGND VGND VPWR VPWR _04940_
+ sky130_fd_sc_hd__mux2_1
X_10086_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__buf_2
Xhold6 rvsingle.dp.rf.rf\[25\]\[20\] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10988_ _04770_ net709 _05419_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12727_ clknet_leaf_6_clk _00185_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12658_ clknet_leaf_41_clk _00116_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11609_ _04972_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12589_ clknet_leaf_44_clk _00047_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_10_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold406 rvsingle.dp.rf.rf\[2\]\[7\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 rvsingle.dp.rf.rf\[26\]\[15\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 rvsingle.dp.rf.rf\[0\]\[16\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold439 rvsingle.dp.rf.rf\[5\]\[19\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _03697_ _01085_ _01837_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__a21oi_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _03666_ _03671_ _02527_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nand3_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07702_ _01125_ rvsingle.dp.rf.rf\[4\]\[5\] _01519_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__o21bai_1
X_08682_ _01780_ rvsingle.dp.rf.rf\[24\]\[14\] VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07633_ rvsingle.dp.rf.rf\[31\]\[4\] _02288_ _02553_ VGND VGND VPWR VPWR _02554_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07564_ _01091_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09303_ _01685_ _04212_ _04217_ _04218_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__a2bb2oi_4
X_06515_ _01306_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__buf_6
XFILLER_0_158_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07495_ rvsingle.dp.rf.rf\[1\]\[6\] _01613_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__and2b_1
XFILLER_0_146_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06446_ rvsingle.dp.rf.rf\[8\]\[28\] rvsingle.dp.rf.rf\[9\]\[28\] rvsingle.dp.rf.rf\[10\]\[28\]
+ rvsingle.dp.rf.rf\[11\]\[28\] _01338_ _01303_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09234_ _02751_ _02857_ _04151_ _04152_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_145_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09165_ _01232_ _04084_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__or2_1
X_06377_ _01197_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08116_ _01769_ rvsingle.dp.rf.rf\[28\]\[1\] _01091_ VGND VGND VPWR VPWR _03037_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09096_ _03857_ rvsingle.dp.rf.rf\[3\]\[26\] _03840_ _04015_ VGND VGND VPWR VPWR
+ _04016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08047_ _02163_ rvsingle.dp.rf.rf\[10\]\[1\] VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09998_ _02909_ _02799_ _02910_ ReadData[15] _04715_ VGND VGND VPWR VPWR _04810_
+ sky130_fd_sc_hd__o311a_1
X_08949_ _01257_ rvsingle.dp.rf.rf\[8\]\[25\] _03869_ _01856_ VGND VGND VPWR VPWR
+ _03870_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_99_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_68_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
X_11960_ _05946_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10911_ _04770_ rvsingle.dp.rf.rf\[18\]\[6\] _05373_ VGND VGND VPWR VPWR _05380_
+ sky130_fd_sc_hd__mux2_1
X_11891_ _04773_ net487 _05902_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10842_ _04915_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10773_ _04828_ rvsingle.dp.rf.rf\[20\]\[18\] _05285_ VGND VGND VPWR VPWR _05294_
+ sky130_fd_sc_hd__mux2_1
X_12512_ clknet_leaf_119_clk _00996_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12443_ clknet_leaf_136_clk _00927_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12374_ clknet_leaf_25_clk _00858_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11325_ _05606_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__buf_6
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11256_ _05318_ rvsingle.dp.rf.rf\[15\]\[1\] _05569_ VGND VGND VPWR VPWR _05570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10207_ _04966_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__clkbuf_8
X_11187_ _04754_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__buf_2
X_10138_ _04931_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_59_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
X_10069_ _04870_ net759 _04847_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06300_ _01222_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__buf_4
X_07280_ rvsingle.dp.rf.rf\[1\]\[16\] _01296_ _01309_ _02200_ VGND VGND VPWR VPWR
+ _02201_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_73_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06231_ _01115_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06162_ Instr[20] VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold203 rvsingle.dp.rf.rf\[3\]\[4\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 rvsingle.dp.rf.rf\[9\]\[26\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 rvsingle.dp.rf.rf\[4\]\[27\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold236 rvsingle.dp.rf.rf\[25\]\[28\] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold247 rvsingle.dp.rf.rf\[8\]\[30\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 rvsingle.dp.rf.rf\[30\]\[30\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _04397_ _04743_ _04744_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__o2bb2a_4
Xhold269 rvsingle.dp.rf.rf\[23\]\[9\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ PC[28] _04663_ PC[29] VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__a21oi_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _03721_ _01689_ _02273_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__a211o_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _04590_ PC[23] VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__nand2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ rvsingle.dp.rf.rf\[8\]\[22\] rvsingle.dp.rf.rf\[9\]\[22\] rvsingle.dp.rf.rf\[10\]\[22\]
+ rvsingle.dp.rf.rf\[11\]\[22\] _01242_ _01434_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__mux4_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _03651_ _03652_ _03654_ _02483_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__o211ai_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _01247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08665_ _01316_ _03579_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__nand3_2
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ rvsingle.dp.rf.rf\[13\]\[4\] _01440_ _01436_ _02536_ VGND VGND VPWR VPWR
+ _02537_ sky130_fd_sc_hd__o211ai_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ rvsingle.dp.rf.rf\[11\]\[12\] _01492_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__or2b_1
XFILLER_0_76_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07547_ _02465_ _02466_ _02467_ _02377_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_165_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07478_ _01860_ rvsingle.dp.rf.rf\[21\]\[6\] _02398_ VGND VGND VPWR VPWR _02399_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09217_ _04135_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__buf_8
XFILLER_0_133_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06429_ _01350_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09148_ _01226_ _04067_ _01210_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09079_ _01943_ rvsingle.dp.rf.rf\[15\]\[26\] _01200_ _03998_ VGND VGND VPWR VPWR
+ _03999_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ _05314_ _05487_ _05488_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12090_ _06014_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__clkbuf_1
Xhold770 rvsingle.dp.rf.rf\[24\]\[22\] VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 rvsingle.dp.rf.rf\[18\]\[24\] VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _05453_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
Xhold792 rvsingle.dp.rf.rf\[8\]\[7\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12992_ clknet_leaf_115_clk _00450_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11943_ _05935_ _05899_ _05936_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _04720_ _04728_ _05830_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__and3_2
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10825_ _04764_ _05316_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__and2_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10756_ _05284_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10687_ _04790_ rvsingle.dp.rf.rf\[21\]\[11\] _05246_ VGND VGND VPWR VPWR _05247_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12426_ clknet_leaf_82_clk _00910_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12357_ _06130_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11308_ _05407_ net508 _05591_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12288_ _04903_ net474 _06073_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__mux2_1
X_11239_ _05307_ net621 _05552_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__mux2_1
X_06780_ _01230_ _01686_ _01700_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_171_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08450_ _01468_ rvsingle.dp.rf.rf\[14\]\[9\] _01198_ VGND VGND VPWR VPWR _03371_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07401_ rvsingle.dp.rf.rf\[13\]\[7\] _01618_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__and2b_1
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08381_ rvsingle.dp.rf.rf\[28\]\[8\] rvsingle.dp.rf.rf\[29\]\[8\] rvsingle.dp.rf.rf\[30\]\[8\]
+ rvsingle.dp.rf.rf\[31\]\[8\] _01730_ _01953_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07332_ rvsingle.dp.rf.rf\[11\]\[16\] _01488_ _02252_ VGND VGND VPWR VPWR _02253_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07263_ _02182_ _02183_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_143_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09002_ _03919_ _01310_ _01915_ _03921_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__a211o_1
X_06214_ _01137_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07194_ rvsingle.dp.rf.rf\[17\]\[17\] _01499_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__and2b_1
XFILLER_0_171_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06145_ Instr[3] Instr[2] _01068_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__nor3_1
XFILLER_0_131_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_997 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09904_ _04719_ _04729_ _04730_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _04617_ PC[27] VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__xnor2_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _04367_ _04599_ _04603_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[21\] sky130_fd_sc_hd__o21ai_1
X_06978_ rvsingle.dp.rf.rf\[20\]\[22\] rvsingle.dp.rf.rf\[21\]\[22\] rvsingle.dp.rf.rf\[22\]\[22\]
+ rvsingle.dp.rf.rf\[23\]\[22\] _01417_ _01301_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__mux4_1
X_08717_ rvsingle.dp.rf.rf\[5\]\[14\] _03258_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__and2b_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _04539_ _04540_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _03467_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__inv_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08579_ _02303_ rvsingle.dp.rf.rf\[27\]\[12\] _01199_ _03499_ VGND VGND VPWR VPWR
+ _03500_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10610_ _05203_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11590_ _05755_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10541_ _04790_ net767 _05152_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13260_ clknet_leaf_93_clk _00718_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10472_ _04818_ net237 _05110_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12211_ reset VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__buf_4
X_13191_ clknet_leaf_101_clk _00649_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12142_ _06041_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12073_ _05639_ net247 _05994_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__mux2_1
X_11024_ _05300_ rvsingle.dp.rf.rf\[31\]\[22\] _05443_ VGND VGND VPWR VPWR _05445_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ clknet_leaf_40_clk _00433_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _05927_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11857_ _05890_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10808_ _05097_ _04726_ _05058_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__and3_2
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11788_ _04876_ net660 _05845_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10739_ _04747_ net790 _05274_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12409_ clknet_leaf_32_clk _00893_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13389_ clknet_leaf_46_clk _00817_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07950_ rvsingle.dp.rf.rf\[7\]\[0\] _01842_ _02870_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__o21ai_1
X_06901_ _01230_ _01821_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__nor2_1
X_07881_ _02801_ _02375_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09620_ Instr[29] PC[9] VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__and2_1
X_06832_ _01752_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09551_ PC[3] _02748_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__nor2_1
X_06763_ _01592_ _01641_ _01683_ _01481_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__nand4_2
XFILLER_0_78_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08502_ _01779_ rvsingle.dp.rf.rf\[20\]\[13\] _01610_ VGND VGND VPWR VPWR _03423_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06694_ _01614_ rvsingle.dp.rf.rf\[12\]\[20\] VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__nor2_1
X_09482_ _01154_ _01774_ _01802_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__and3_2
XFILLER_0_53_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08433_ rvsingle.dp.rf.rf\[17\]\[9\] _01607_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08364_ _01328_ rvsingle.dp.rf.rf\[6\]\[8\] VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07315_ _01768_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08295_ _03208_ _03210_ _02527_ _03215_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_15_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07246_ _01722_ _02160_ _01478_ _02166_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_116_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07177_ _02066_ _02068_ _02081_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09818_ _04590_ PC[26] VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__nand2_1
X_09749_ PC[19] _04577_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ clknet_leaf_34_clk _00218_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _05295_ rvsingle.dp.rf.rf\[10\]\[19\] _05806_ VGND VGND VPWR VPWR _05815_
+ sky130_fd_sc_hd__mux2_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12691_ clknet_leaf_28_clk _00149_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11642_ _04818_ _04973_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11573_ _04802_ _04973_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13312_ clknet_leaf_133_clk _00770_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10524_ _05113_ _05114_ _05115_ _05061_ _04754_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__o311a_1
XFILLER_0_162_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13243_ clknet_leaf_10_clk _00701_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10455_ _04879_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13174_ clknet_leaf_62_clk _00632_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10386_ _04786_ rvsingle.dp.rf.rf\[25\]\[10\] _05071_ VGND VGND VPWR VPWR _05075_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12125_ _04845_ net791 _06031_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12056_ _04845_ net666 _05994_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11007_ _05435_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12958_ clknet_leaf_150_clk _00416_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11909_ _05918_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12889_ clknet_leaf_8_clk _00347_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_270 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_281 _02314_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_292 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07100_ _02017_ _02018_ _01132_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_160_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08080_ _01797_ rvsingle.dp.rf.rf\[0\]\[1\] _03000_ _01667_ VGND VGND VPWR VPWR _03001_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07031_ rvsingle.dp.rf.rf\[1\]\[19\] _01441_ _01689_ _01951_ VGND VGND VPWR VPWR
+ _01952_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08982_ _01463_ rvsingle.dp.rf.rf\[2\]\[25\] VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__or2_1
X_07933_ _01188_ _02682_ _02695_ _01247_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__o211a_1
X_07864_ _02779_ _02784_ _01505_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__nand3_1
XFILLER_0_74_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09603_ _04363_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__buf_2
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06815_ _01720_ _01724_ _01188_ _01735_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__o211ai_2
X_07795_ rvsingle.dp.rf.rf\[5\]\[3\] _01779_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__and2b_1
X_09534_ _04305_ _04306_ VGND VGND VPWR VPWR DataAdr[24] sky130_fd_sc_hd__nand2_8
XFILLER_0_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06746_ _01091_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09465_ _01094_ net825 _03044_ _01058_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__o211ai_1
X_06677_ rvsingle.dp.rf.rf\[9\]\[20\] _01097_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08416_ rvsingle.dp.rf.rf\[7\]\[9\] _01492_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__or2b_1
XFILLER_0_164_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09396_ _02377_ _02374_ _02468_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08347_ _03264_ _03267_ _01505_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_129_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08278_ _01105_ _03195_ _03196_ _02483_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07229_ _01962_ _01100_ _02126_ _02149_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_81_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10240_ _04786_ rvsingle.dp.rf.rf\[27\]\[10\] _04989_ VGND VGND VPWR VPWR _04993_
+ sky130_fd_sc_hd__mux2_1
X_10171_ _04948_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12812_ clknet_leaf_50_clk _00270_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ clknet_leaf_98_clk _00201_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12674_ clknet_leaf_128_clk _00132_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11625_ _05777_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11556_ net125 _05731_ _05736_ _05737_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10507_ _04915_ _04965_ _04917_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11487_ _05683_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__buf_6
X_13226_ clknet_leaf_102_clk _00684_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10438_ _04736_ net771 _05103_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ clknet_leaf_115_clk _00615_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10369_ _05066_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__clkbuf_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _04801_ net554 _06019_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ clknet_leaf_119_clk _00546_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12039_ _05976_ net168 _05119_ _05146_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_06600_ _01518_ rvsingle.dp.rf.rf\[20\]\[21\] _01520_ VGND VGND VPWR VPWR _01521_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_88_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07580_ rvsingle.dp.rf.rf\[13\]\[4\] _01508_ _02395_ VGND VGND VPWR VPWR _02501_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06531_ _01451_ _01351_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__nor2_8
XFILLER_0_76_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09250_ _01927_ _01929_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06462_ _01383_ rvsingle.dp.rf.rf\[30\]\[28\] VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08201_ _03118_ _03119_ _02543_ _03121_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_118_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06393_ Instr[19] VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__inv_6
X_09181_ rvsingle.dp.rf.rf\[8\]\[31\] rvsingle.dp.rf.rf\[9\]\[31\] rvsingle.dp.rf.rf\[10\]\[31\]
+ rvsingle.dp.rf.rf\[11\]\[31\] _01100_ _01120_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08132_ _02967_ _03049_ _03047_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08063_ _01191_ rvsingle.dp.rf.rf\[18\]\[1\] VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07014_ _01230_ _01934_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08965_ _01194_ rvsingle.dp.rf.rf\[18\]\[25\] VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__or2_1
X_07916_ _01462_ rvsingle.dp.rf.rf\[24\]\[2\] _01299_ VGND VGND VPWR VPWR _02837_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08896_ _03815_ _03816_ _01445_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__mux2_1
X_07847_ _01675_ rvsingle.dp.rf.rf\[4\]\[2\] VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__nor2_1
X_07778_ _01097_ rvsingle.dp.rf.rf\[8\]\[3\] VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09517_ _04394_ VGND VGND VPWR VPWR WriteData[1] sky130_fd_sc_hd__clkbuf_4
X_06729_ _01135_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__buf_6
XFILLER_0_67_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _03056_ _02576_ _02667_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09379_ net821 _03141_ _03230_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__o21ai_2
X_11410_ _05653_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12390_ clknet_leaf_121_clk _00874_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11341_ _05615_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11272_ _05428_ net501 _05569_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13011_ clknet_leaf_29_clk _00469_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10223_ _04917_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__clkbuf_4
X_10154_ _04939_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
X_10085_ _04365_ _04883_ _04884_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__o21bai_4
Xhold7 rvsingle.dp.rf.rf\[27\]\[0\] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10987_ _05424_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12726_ clknet_leaf_32_clk _00184_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12657_ clknet_leaf_49_clk _00115_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11608_ _05765_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12588_ clknet_leaf_49_clk _00046_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11539_ _04976_ _04975_ _05149_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__or3_2
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold407 rvsingle.dp.rf.rf\[15\]\[30\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 rvsingle.dp.rf.rf\[26\]\[18\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold429 rvsingle.dp.rf.rf\[16\]\[29\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13209_ clknet_leaf_15_clk _00667_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _01531_ _03667_ _03668_ _01131_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__o311ai_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07701_ _02379_ rvsingle.dp.rf.rf\[7\]\[5\] _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__o21a_1
X_08681_ _03598_ _03599_ _03601_ _01617_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_135_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07632_ _01725_ rvsingle.dp.rf.rf\[30\]\[4\] _01198_ VGND VGND VPWR VPWR _02553_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07563_ _02477_ _02479_ _02480_ _02482_ _02483_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09302_ _04167_ _01742_ _04125_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06514_ rvsingle.dp.rf.rf\[16\]\[21\] rvsingle.dp.rf.rf\[17\]\[21\] rvsingle.dp.rf.rf\[18\]\[21\]
+ rvsingle.dp.rf.rf\[19\]\[21\] _01432_ _01434_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07494_ _02117_ rvsingle.dp.rf.rf\[0\]\[6\] VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09233_ _02851_ _02803_ _02856_ _02751_ _02861_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__o2111ai_4
X_06445_ _01363_ _01365_ _01210_ _01366_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_61_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09164_ rvsingle.dp.rf.rf\[24\]\[31\] rvsingle.dp.rf.rf\[25\]\[31\] rvsingle.dp.rf.rf\[26\]\[31\]
+ rvsingle.dp.rf.rf\[27\]\[31\] _01196_ _01203_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06376_ _01297_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08115_ rvsingle.dp.rf.rf\[29\]\[1\] _01544_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__and2b_1
X_09095_ _01126_ rvsingle.dp.rf.rf\[2\]\[26\] VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_783 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08046_ _02907_ _02963_ _02966_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_114_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09997_ _04809_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__clkbuf_1
X_08948_ rvsingle.dp.rf.rf\[9\]\[25\] _01126_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__or2b_1
X_08879_ _02236_ _03795_ _03799_ _01157_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__o211ai_1
X_10910_ _05379_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__clkbuf_1
X_11890_ _05908_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10841_ _05316_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10772_ _05293_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12511_ clknet_leaf_13_clk _00995_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12442_ clknet_leaf_4_clk _00926_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12373_ clknet_leaf_60_clk _00857_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11324_ _05565_ _04738_ _04739_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__or3b_4
X_11255_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__buf_6
X_10206_ _04720_ _04966_ _04967_ _04968_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__and4_2
X_11186_ _05530_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10137_ _04736_ rvsingle.dp.rf.rf\[28\]\[1\] _04930_ VGND VGND VPWR VPWR _04931_
+ sky130_fd_sc_hd__mux2_1
X_10068_ _04869_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12709_ clknet_leaf_110_clk _00167_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06230_ _01153_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06161_ _01084_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold204 rvsingle.dp.rf.rf\[19\]\[3\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 rvsingle.dp.rf.rf\[5\]\[27\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 rvsingle.dp.rf.rf\[30\]\[23\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold237 rvsingle.dp.rf.rf\[24\]\[16\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold248 rvsingle.dp.rf.rf\[11\]\[0\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _04364_ _04141_ _04732_ DataAdr[2] VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__o31a_1
Xhold259 rvsingle.dp.rf.rf\[10\]\[24\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ PC[27] PC[28] _04660_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__and3_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _02929_ rvsingle.dp.rf.rf\[3\]\[15\] _01727_ _03722_ VGND VGND VPWR VPWR
+ _03723_ sky130_fd_sc_hd__o211a_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _04617_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__buf_2
X_06994_ _01694_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__clkbuf_8
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _01878_ rvsingle.dp.rf.rf\[16\]\[15\] _03653_ _02395_ VGND VGND VPWR VPWR
+ _03654_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _03580_ _01445_ _01699_ _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_96_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _01419_ rvsingle.dp.rf.rf\[12\]\[4\] VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _03514_ _03515_ _01131_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_165_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07546_ _01065_ _01074_ _01870_ _02319_ _02372_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__o221a_1
XFILLER_0_165_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07477_ _01544_ rvsingle.dp.rf.rf\[20\]\[6\] _01610_ VGND VGND VPWR VPWR _02398_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09216_ _04121_ _04122_ _04117_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__o21a_4
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06428_ _01349_ Instr[17] _01215_ Instr[19] VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09147_ rvsingle.dp.rf.rf\[14\]\[31\] rvsingle.dp.rf.rf\[15\]\[31\] _01196_ VGND
+ VGND VPWR VPWR _04067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06359_ _01099_ rvsingle.dp.rf.rf\[24\]\[29\] VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09078_ _01432_ rvsingle.dp.rf.rf\[14\]\[26\] VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08029_ rvsingle.dp.rf.rf\[0\]\[0\] _02440_ _01454_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__o21bai_1
Xhold760 rvsingle.dp.rf.rf\[30\]\[18\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 rvsingle.dp.rf.rf\[24\]\[1\] VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold782 rvsingle.dp.rf.rf\[20\]\[10\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _05187_ net426 _05443_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__mux2_1
Xhold793 rvsingle.dp.rf.rf\[16\]\[21\] VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12991_ clknet_leaf_2_clk _00449_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11942_ _05769_ _05770_ _05899_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__o21ai_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _05898_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__inv_2
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10824_ _05085_ _05326_ _05325_ net193 VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10755_ _04786_ net782 _05274_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10686_ _05234_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__buf_6
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12425_ clknet_leaf_94_clk _00909_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12356_ _04897_ net261 _06121_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11307_ _05596_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__clkbuf_1
X_12287_ _04898_ _05145_ _05832_ _06092_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11238_ _05558_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__clkbuf_1
X_11169_ _05359_ net351 _05511_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07400_ _01862_ rvsingle.dp.rf.rf\[12\]\[7\] VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08380_ _01200_ _03298_ _03300_ _01694_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_19_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07331_ _01562_ rvsingle.dp.rf.rf\[10\]\[16\] _01620_ VGND VGND VPWR VPWR _02252_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07262_ _02181_ _02151_ _02153_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__nand3_1
X_09001_ _01943_ rvsingle.dp.rf.rf\[19\]\[27\] _01451_ _03920_ VGND VGND VPWR VPWR
+ _03921_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06213_ _01136_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__clkbuf_8
X_07193_ _01603_ rvsingle.dp.rf.rf\[16\]\[17\] _02031_ VGND VGND VPWR VPWR _02114_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_26_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06144_ Instr[4] Instr[1] Instr[0] Instr[5] VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_130_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09903_ net35 _04729_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__nor2_1
Xwire5 _02911_ VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__buf_1
XFILLER_0_10_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09834_ _04618_ PC[26] _04650_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__o21bai_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _04398_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__nand2_1
X_06977_ _01591_ _01580_ _01897_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__and3_1
X_08716_ _01567_ rvsingle.dp.rf.rf\[4\]\[14\] VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ PC[14] _04529_ _04531_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__a21oi_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08647_ _01316_ _03473_ _03480_ _01452_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__a31o_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _01462_ rvsingle.dp.rf.rf\[26\]\[12\] VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07529_ _01327_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__buf_8
XFILLER_0_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10540_ net50 _05155_ _05164_ _05157_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10471_ _05122_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12210_ _05898_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13190_ clknet_leaf_111_clk _00648_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12141_ _05716_ net219 _06031_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12072_ _06003_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__clkbuf_1
Xhold590 rvsingle.dp.rf.rf\[14\]\[4\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11023_ _05444_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__clkbuf_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ clknet_leaf_52_clk _00432_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _05757_ rvsingle.dp.rf.rf\[6\]\[23\] _05924_ VGND VGND VPWR VPWR _05927_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _04869_ net477 _05885_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__mux2_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10807_ _04718_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11787_ _05837_ net190 _05760_ _05841_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10738_ _05275_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10669_ _05237_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12408_ clknet_leaf_34_clk _00892_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13388_ clknet_leaf_51_clk _00816_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12339_ _06098_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__buf_8
X_06900_ rvsingle.dp.rf.rf\[16\]\[23\] rvsingle.dp.rf.rf\[17\]\[23\] rvsingle.dp.rf.rf\[18\]\[23\]
+ rvsingle.dp.rf.rf\[19\]\[23\] _01329_ _01456_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__mux4_1
X_07880_ _01512_ net825 _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__o21a_2
XFILLER_0_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06831_ Instr[20] VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__buf_4
X_09550_ _04397_ PC[3] VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__xnor2_2
X_06762_ _01664_ _01681_ _01682_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__nand3_4
XFILLER_0_78_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08501_ _01097_ rvsingle.dp.rf.rf\[18\]\[13\] _01654_ _03421_ VGND VGND VPWR VPWR
+ _03422_ sky130_fd_sc_hd__o211a_1
X_09481_ _04381_ VGND VGND VPWR VPWR WriteData[24] sky130_fd_sc_hd__clkbuf_4
X_06693_ _01613_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08432_ _02030_ rvsingle.dp.rf.rf\[16\]\[9\] _01104_ VGND VGND VPWR VPWR _03353_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_53_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08363_ rvsingle.dp.rf.rf\[4\]\[8\] rvsingle.dp.rf.rf\[5\]\[8\] _01420_ VGND VGND
+ VPWR VPWR _03284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07314_ rvsingle.dp.rf.rf\[4\]\[16\] rvsingle.dp.rf.rf\[5\]\[16\] _01666_ VGND VGND
+ VPWR VPWR _02235_ sky130_fd_sc_hd__mux2_1
X_08294_ _01605_ _03211_ _03212_ _01511_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_15_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07245_ _02161_ _01437_ _01702_ _02165_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07176_ _02088_ _01450_ _02096_ _01452_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__a31o_2
XFILLER_0_41_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09817_ _04636_ _04648_ _04649_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__a21oi_1
X_09748_ _04568_ _04572_ _04586_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__a21o_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _04454_ _04455_ _04524_ _04459_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__o211ai_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _05814_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__clkbuf_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12690_ clknet_leaf_27_clk _00148_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11641_ _05471_ _05749_ _05779_ net202 VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_139_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11572_ _05167_ _05746_ _05731_ net143 VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_25_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13311_ clknet_leaf_135_clk _00769_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10523_ _05152_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13242_ clknet_leaf_22_clk _00700_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_10454_ _05112_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13173_ clknet_leaf_17_clk _00631_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10385_ _05074_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__clkbuf_1
X_12124_ _06032_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__clkbuf_1
X_12055_ _05976_ net161 _05149_ _05513_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__o2bb2ai_1
X_11006_ _05391_ rvsingle.dp.rf.rf\[31\]\[14\] _05431_ VGND VGND VPWR VPWR _05435_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ clknet_leaf_142_clk _00415_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ _04813_ net561 _05913_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_260 _01531_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12888_ clknet_leaf_32_clk _00346_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_271 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_282 _02314_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_293 _05271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11839_ _05476_ net562 _05874_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07030_ _01707_ rvsingle.dp.rf.rf\[0\]\[19\] VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08981_ rvsingle.dp.rf.rf\[0\]\[25\] rvsingle.dp.rf.rf\[1\]\[25\] _01336_ VGND VGND
+ VPWR VPWR _03901_ sky130_fd_sc_hd__mux2_1
X_07932_ _02852_ _01584_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__nand2_1
X_07863_ _01552_ _02780_ _02781_ _02329_ _02783_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__o311ai_2
X_06814_ _01703_ _01729_ _01734_ _01478_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__o211ai_1
X_09602_ _04139_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__buf_2
X_07794_ _01125_ rvsingle.dp.rf.rf\[4\]\[3\] VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__nor2_1
X_09533_ _04210_ VGND VGND VPWR VPWR DataAdr[22] sky130_fd_sc_hd__clkinv_4
XFILLER_0_79_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06745_ _01148_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09464_ PC[1] _03045_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06676_ _01595_ rvsingle.dp.rf.rf\[8\]\[20\] _01596_ VGND VGND VPWR VPWR _01597_
+ sky130_fd_sc_hd__o21bai_1
X_08415_ rvsingle.dp.rf.rf\[5\]\[9\] _01743_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09395_ _04308_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08346_ _03265_ _03266_ _02351_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08277_ _01268_ rvsingle.dp.rf.rf\[18\]\[10\] _02059_ _03197_ VGND VGND VPWR VPWR
+ _03198_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07228_ _01593_ _02137_ _02148_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__nand3_4
XFILLER_0_131_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07159_ _01915_ _02075_ _02077_ _02079_ _01222_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__o221ai_4
X_10170_ _04824_ net755 _04941_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12811_ clknet_leaf_86_clk _00269_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[16\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ clknet_leaf_113_clk _00200_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ clknet_leaf_140_clk _00131_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11624_ _05728_ net483 _05775_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11555_ _05146_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10506_ _05140_ _05098_ _05141_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11486_ _05694_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13225_ clknet_leaf_127_clk _00683_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10437_ _05102_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__buf_8
XFILLER_0_0_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13156_ clknet_leaf_109_clk _00614_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10368_ _04736_ net370 _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__mux2_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _06023_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__clkbuf_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ clknet_leaf_2_clk _00545_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10299_ _04760_ net416 _05022_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__mux2_1
X_12038_ _05987_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06530_ _01244_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__buf_8
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06461_ _01382_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_919 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08200_ rvsingle.dp.rf.rf\[9\]\[11\] _02303_ _01308_ _03120_ VGND VGND VPWR VPWR
+ _03121_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09180_ rvsingle.dp.rf.rf\[12\]\[31\] rvsingle.dp.rf.rf\[13\]\[31\] rvsingle.dp.rf.rf\[14\]\[31\]
+ rvsingle.dp.rf.rf\[15\]\[31\] _01100_ _01120_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06392_ _01210_ _01305_ _01313_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08131_ _03050_ _03051_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08062_ rvsingle.dp.rf.rf\[16\]\[1\] rvsingle.dp.rf.rf\[17\]\[1\] _01241_ VGND VGND
+ VPWR VPWR _02983_ sky130_fd_sc_hd__mux2_1
X_07013_ rvsingle.dp.rf.rf\[16\]\[19\] rvsingle.dp.rf.rf\[17\]\[19\] rvsingle.dp.rf.rf\[18\]\[19\]
+ rvsingle.dp.rf.rf\[19\]\[19\] _01329_ _01456_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08964_ rvsingle.dp.rf.rf\[16\]\[25\] rvsingle.dp.rf.rf\[17\]\[25\] _01194_ VGND
+ VGND VPWR VPWR _03884_ sky130_fd_sc_hd__mux2_1
X_07915_ _02543_ _02833_ _02835_ _01215_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__a31o_1
X_08895_ rvsingle.dp.rf.rf\[4\]\[24\] rvsingle.dp.rf.rf\[5\]\[24\] rvsingle.dp.rf.rf\[6\]\[24\]
+ rvsingle.dp.rf.rf\[7\]\[24\] _01726_ _01728_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__mux4_1
X_07846_ _01567_ rvsingle.dp.rf.rf\[2\]\[2\] _02031_ _02766_ VGND VGND VPWR VPWR _02767_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07777_ Instr[10] _01078_ _02697_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_79_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06728_ rvsingle.dp.rf.rf\[31\]\[20\] _01646_ _01648_ VGND VGND VPWR VPWR _01649_
+ sky130_fd_sc_hd__o21ai_1
X_09516_ _04377_ _03019_ _03042_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__and3_2
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _04351_ _04136_ _04352_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_164_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06659_ _01171_ _01176_ net822 VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__o21ai_4
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09378_ DataAdr[18] VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08329_ rvsingle.dp.rf.rf\[7\]\[8\] _01487_ _01523_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11340_ _05330_ net708 _05607_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11271_ _05577_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__clkbuf_1
X_13010_ clknet_leaf_57_clk _00468_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10222_ _04915_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10153_ _04782_ net600 _04930_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__mux2_1
X_10084_ _04425_ _04665_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__nor2_1
Xhold8 rvsingle.dp.rf.rf\[24\]\[9\] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10986_ _04765_ rvsingle.dp.rf.rf\[31\]\[5\] _05419_ VGND VGND VPWR VPWR _05424_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12725_ clknet_leaf_58_clk _00183_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12656_ clknet_leaf_72_clk _00114_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11607_ _05716_ net255 _05729_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12587_ clknet_leaf_87_clk _00045_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11538_ _04735_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__buf_2
XFILLER_0_64_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold408 rvsingle.dp.rf.rf\[17\]\[28\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold419 rvsingle.dp.rf.rf\[29\]\[8\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _05322_ net253 _05684_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13208_ clknet_leaf_22_clk _00666_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13139_ clknet_leaf_28_clk _00597_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _01566_ rvsingle.dp.rf.rf\[6\]\[5\] _01258_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__o21a_1
X_08680_ rvsingle.dp.rf.rf\[29\]\[14\] _02481_ _01496_ _03600_ VGND VGND VPWR VPWR
+ _03601_ sky130_fd_sc_hd__o211ai_1
X_07631_ rvsingle.dp.rf.rf\[29\]\[4\] _02275_ _01436_ _02551_ VGND VGND VPWR VPWR
+ _02552_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07562_ _01599_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09301_ _04215_ _04216_ _03767_ _01742_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__a31o_1
X_06513_ _01433_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07493_ _02404_ _02407_ _01505_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_146_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09232_ _03047_ _03052_ _02967_ _03049_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__a2bb2oi_4
X_06444_ rvsingle.dp.rf.rf\[4\]\[28\] rvsingle.dp.rf.rf\[5\]\[28\] rvsingle.dp.rf.rf\[6\]\[28\]
+ rvsingle.dp.rf.rf\[7\]\[28\] _01338_ _01202_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09163_ _01298_ rvsingle.dp.rf.rf\[31\]\[31\] _01226_ _04082_ VGND VGND VPWR VPWR
+ _04083_ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06375_ _01296_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08114_ _01259_ _03031_ _03032_ _01599_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__o311ai_1
X_09094_ rvsingle.dp.rf.rf\[0\]\[26\] rvsingle.dp.rf.rf\[1\]\[26\] _01269_ VGND VGND
+ VPWR VPWR _04014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08045_ _02964_ _02965_ _01183_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__nand3_2
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09996_ _04808_ net602 _04791_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08947_ rvsingle.dp.rf.rf\[11\]\[25\] _03857_ _03840_ VGND VGND VPWR VPWR _03868_
+ sky130_fd_sc_hd__o21ai_1
X_08878_ _03796_ _01543_ _01632_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07829_ _02749_ _02746_ _01485_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10840_ _05335_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10771_ _04824_ net485 _05285_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_145_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_145_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12510_ clknet_leaf_135_clk _00994_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12441_ clknet_leaf_7_clk _00925_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12372_ clknet_leaf_21_clk _00856_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11323_ _05314_ _05604_ _05605_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11254_ _05417_ _05565_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or2_2
X_10205_ _04739_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__buf_2
X_11185_ _05322_ net805 _05528_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10136_ _04929_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__buf_8
X_10067_ _04868_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_136_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_136_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10969_ net56 VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12708_ clknet_leaf_124_clk _00166_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12639_ clknet_leaf_2_clk _00097_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06160_ _01083_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_170_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold205 rvsingle.dp.rf.rf\[1\]\[20\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold216 rvsingle.dp.rf.rf\[24\]\[28\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 rvsingle.dp.rf.rf\[2\]\[15\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold238 rvsingle.dp.rf.rf\[1\]\[23\] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 rvsingle.dp.rf.rf\[6\]\[24\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _04678_ _04452_ _04680_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[28\] sky130_fd_sc_hd__o21ai_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _01240_ rvsingle.dp.rf.rf\[2\]\[15\] VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__or2_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _01222_ _01907_ _01913_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__o21ai_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _04590_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__clkbuf_4
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ rvsingle.dp.rf.rf\[17\]\[15\] _01877_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__or2b_1
X_08663_ _03581_ _01716_ _01460_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07614_ rvsingle.dp.rf.rf\[8\]\[4\] rvsingle.dp.rf.rf\[9\]\[4\] rvsingle.dp.rf.rf\[10\]\[4\]
+ rvsingle.dp.rf.rf\[11\]\[4\] _01416_ _01708_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__mux4_1
X_08594_ rvsingle.dp.rf.rf\[9\]\[12\] _03258_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__and2b_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07545_ _02301_ _02314_ _01188_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_127_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_127_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07476_ rvsingle.dp.rf.rf\[23\]\[6\] _01594_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__and2b_1
XFILLER_0_147_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09215_ _01250_ _04063_ _04116_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__nand3_1
X_06427_ _01190_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09146_ rvsingle.dp.rf.rf\[13\]\[31\] _01298_ _01311_ _04065_ VGND VGND VPWR VPWR
+ _04066_ sky130_fd_sc_hd__o211a_1
X_06358_ rvsingle.dp.rf.rf\[27\]\[29\] _01090_ _01280_ VGND VGND VPWR VPWR _01281_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09077_ rvsingle.dp.rf.rf\[12\]\[26\] rvsingle.dp.rf.rf\[13\]\[26\] _01193_ VGND
+ VGND VPWR VPWR _03997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06289_ rvsingle.dp.rf.rf\[4\]\[30\] rvsingle.dp.rf.rf\[5\]\[30\] rvsingle.dp.rf.rf\[6\]\[30\]
+ rvsingle.dp.rf.rf\[7\]\[30\] _01196_ _01203_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08028_ _01444_ _02941_ _02943_ _01215_ _02948_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__o311ai_1
Xhold750 rvsingle.dp.rf.rf\[21\]\[27\] VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 rvsingle.dp.rf.rf\[14\]\[15\] VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 rvsingle.dp.rf.rf\[31\]\[24\] VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 rvsingle.dp.rf.rf\[21\]\[2\] VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold794 rvsingle.dp.rf.rf\[20\]\[20\] VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__dlygate4sd3_1
X_09979_ _04793_ _04513_ _04364_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__mux2_4
X_12990_ clknet_leaf_150_clk _00448_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11941_ net43 VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__inv_2
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _05898_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__inv_2
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _04982_ _04983_ _04981_ _04759_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__or4b_2
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_118_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_118_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10754_ _05283_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10685_ _05245_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12424_ clknet_leaf_106_clk _00908_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12355_ _06129_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11306_ _05304_ rvsingle.dp.rf.rf\[15\]\[25\] _05591_ VGND VGND VPWR VPWR _05596_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12286_ _05084_ _05835_ net276 VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__o21a_1
X_11237_ _05407_ net603 _05552_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11168_ _05519_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__clkbuf_1
X_10119_ _04906_ _04729_ _04914_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__o21ai_1
X_11099_ _05359_ net408 _05469_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_109_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_109_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07330_ rvsingle.dp.rf.rf\[9\]\[16\] _01509_ _01543_ VGND VGND VPWR VPWR _02251_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07261_ _02151_ _02153_ _02181_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09000_ _01242_ rvsingle.dp.rf.rf\[18\]\[27\] VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06212_ _01135_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__buf_4
X_07192_ _01512_ _02107_ _02112_ _01526_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06143_ Instr[6] VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09902_ _04721_ _04726_ _04728_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__and3_2
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09833_ _04663_ _04664_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__or2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _04600_ _04601_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__xor2_1
X_06976_ _01869_ _01870_ _01592_ _01896_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__nand4_2
X_08715_ _01531_ _03632_ _03633_ _02351_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__o311ai_1
X_09695_ _04537_ _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08646_ _03562_ _03564_ _03497_ _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__o2bb2ai_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ rvsingle.dp.rf.rf\[24\]\[12\] rvsingle.dp.rf.rf\[25\]\[12\] _01691_ VGND
+ VGND VPWR VPWR _03498_ sky130_fd_sc_hd__mux2_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07528_ _02436_ _02439_ _02448_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_18_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07459_ rvsingle.dp.rf.rf\[27\]\[6\] _02379_ _01777_ VGND VGND VPWR VPWR _02380_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10470_ _04814_ rvsingle.dp.rf.rf\[24\]\[15\] _05110_ VGND VGND VPWR VPWR _05122_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09129_ _01117_ _04036_ _04041_ _01147_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_150_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12140_ _06040_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12071_ _05716_ net288 _05994_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold580 rvsingle.dp.rf.rf\[27\]\[25\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold591 rvsingle.dp.rf.rf\[20\]\[26\] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _05400_ rvsingle.dp.rf.rf\[31\]\[21\] _05443_ VGND VGND VPWR VPWR _05444_
+ sky130_fd_sc_hd__mux2_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ clknet_leaf_42_clk _00431_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _05926_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__clkbuf_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _05889_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10806_ _05312_ _05271_ _05313_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__o21ai_1
X_11786_ _05852_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10737_ _04736_ rvsingle.dp.rf.rf\[20\]\[1\] _05274_ VGND VGND VPWR VPWR _05275_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10668_ _04747_ net783 _05235_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12407_ clknet_leaf_6_clk _00891_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13387_ clknet_leaf_87_clk _00815_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10599_ _04760_ net672 _05194_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12338_ _06120_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12269_ _04833_ net439 _06073_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__mux2_1
X_06830_ _01603_ rvsingle.dp.rf.rf\[10\]\[23\] _01605_ _01750_ VGND VGND VPWR VPWR
+ _01751_ sky130_fd_sc_hd__o211ai_1
X_06761_ _01145_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__buf_12
X_08500_ rvsingle.dp.rf.rf\[19\]\[13\] _01381_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__or2b_1
X_09480_ _01154_ _03790_ _03801_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__and3_1
X_06692_ _01095_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08431_ _03346_ _03351_ _01116_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__nand3_1
XFILLER_0_148_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08362_ _03282_ _01584_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07313_ _02217_ _02222_ _01147_ _02233_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_74_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08293_ _01878_ rvsingle.dp.rf.rf\[30\]\[10\] _01520_ _03213_ VGND VGND VPWR VPWR
+ _03214_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07244_ _01440_ rvsingle.dp.rf.rf\[11\]\[17\] _02162_ _02164_ VGND VGND VPWR VPWR
+ _02165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07175_ _01208_ _02090_ _02092_ _02095_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09816_ PC[24] PC[25] _04617_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__o21a_1
X_09747_ _04577_ PC[19] PC[18] _04570_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06959_ _01258_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__buf_6
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _04522_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__nor2_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08629_ _01137_ rvsingle.dp.rf.rf\[28\]\[12\] _03549_ _02485_ VGND VGND VPWR VPWR
+ _03550_ sky130_fd_sc_hd__o211ai_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _05471_ _05748_ _05779_ net126 VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_37_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11571_ _04796_ _04973_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13310_ clknet_leaf_146_clk _00768_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10522_ _05154_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13241_ clknet_leaf_15_clk _00699_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10453_ _04778_ rvsingle.dp.rf.rf\[24\]\[8\] _05110_ VGND VGND VPWR VPWR _05112_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10384_ _04782_ net787 _05071_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13172_ clknet_leaf_56_clk _00630_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12123_ _04839_ net674 _06031_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12054_ _05995_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__clkbuf_1
X_11005_ _05434_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ clknet_leaf_148_clk _00414_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _05917_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__clkbuf_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ clknet_leaf_7_clk _00345_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_250 _01148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_261 _01531_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_272 _01808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _05880_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_283 _04741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_294 _05271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11769_ _05835_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_40_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_960 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08980_ rvsingle.dp.rf.rf\[4\]\[25\] rvsingle.dp.rf.rf\[5\]\[25\] rvsingle.dp.rf.rf\[6\]\[25\]
+ rvsingle.dp.rf.rf\[7\]\[25\] _01330_ _01302_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07931_ _01870_ _02698_ _02746_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07862_ _01862_ rvsingle.dp.rf.rf\[26\]\[2\] _01880_ _02782_ VGND VGND VPWR VPWR
+ _02783_ sky130_fd_sc_hd__o211ai_1
X_09601_ _04452_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__clkbuf_4
X_06813_ _01731_ _01437_ _01721_ _01733_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__a211o_1
X_07793_ _02031_ _02710_ _02711_ _01599_ _02713_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_79_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09532_ _04206_ VGND VGND VPWR VPWR DataAdr[21] sky130_fd_sc_hd__inv_6
X_06744_ rvsingle.dp.rf.rf\[23\]\[20\] VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__inv_2
X_09463_ _04368_ PC[0] _04369_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__and3_1
X_06675_ _01103_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08414_ _01268_ rvsingle.dp.rf.rf\[4\]\[9\] VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09394_ _02464_ _02475_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08345_ rvsingle.dp.rf.rf\[27\]\[8\] _01769_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_31_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08276_ rvsingle.dp.rf.rf\[19\]\[10\] _01492_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07227_ _01634_ _02142_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07158_ _02078_ _01717_ _01722_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07089_ _01990_ _01997_ _02009_ _01593_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__o211ai_4
Xclkbuf_leaf_98_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12810_ clknet_leaf_80_clk _00268_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12741_ clknet_leaf_114_clk _00199_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12672_ clknet_leaf_117_clk _00130_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11623_ _05776_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__clkbuf_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11554_ _04764_ _05732_ _05733_ _05060_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10505_ _04909_ _04913_ _05098_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11485_ _05385_ net653 _05684_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13224_ clknet_leaf_111_clk _00682_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10436_ _04737_ _04919_ _04733_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__or4_4
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13155_ clknet_leaf_118_clk _00613_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10367_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__buf_8
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _04795_ net513 _06019_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__mux2_1
X_10298_ _05025_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__clkbuf_1
X_13086_ clknet_leaf_0_clk _00544_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12037_ _05744_ net218 _05983_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12939_ clknet_leaf_86_clk _00397_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06460_ _01381_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06391_ rvsingle.dp.rf.rf\[1\]\[29\] _01298_ _01311_ _01312_ VGND VGND VPWR VPWR
+ _01313_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08130_ _02473_ _02318_ _03043_ _03046_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08061_ _02974_ _02981_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07012_ _01722_ _01932_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08963_ _01209_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07914_ _01827_ rvsingle.dp.rf.rf\[17\]\[2\] _02834_ VGND VGND VPWR VPWR _02835_
+ sky130_fd_sc_hd__o21ai_1
X_08894_ rvsingle.dp.rf.rf\[0\]\[24\] rvsingle.dp.rf.rf\[1\]\[24\] rvsingle.dp.rf.rf\[2\]\[24\]
+ rvsingle.dp.rf.rf\[3\]\[24\] _01726_ _01728_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__mux4_1
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07845_ rvsingle.dp.rf.rf\[3\]\[2\] _02627_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__or2b_1
XFILLER_0_79_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07776_ _01076_ _01071_ _01062_ _01115_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__a31o_1
X_09515_ _04393_ VGND VGND VPWR VPWR WriteData[2] sky130_fd_sc_hd__clkbuf_4
X_06727_ _01647_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__buf_6
XFILLER_0_66_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ _02665_ _02660_ _04320_ _02666_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__o211a_1
X_06658_ _01482_ _01483_ _01486_ _01578_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__o211a_1
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09377_ _04277_ _04290_ _04292_ VGND VGND VPWR VPWR DataAdr[18] sky130_fd_sc_hd__o21ai_4
XFILLER_0_35_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06589_ rvsingle.dp.rf.rf\[31\]\[21\] _01509_ _01491_ VGND VGND VPWR VPWR _01510_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08328_ _01137_ rvsingle.dp.rf.rf\[6\]\[8\] VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08259_ _02478_ rvsingle.dp.rf.rf\[13\]\[10\] _03179_ VGND VGND VPWR VPWR _03180_
+ sky130_fd_sc_hd__o21ai_2
X_11270_ _05330_ net806 _05569_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10221_ _04965_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10152_ _04938_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__clkbuf_1
X_10083_ _02908_ DataAdr[27] _04882_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__a21oi_1
Xhold9 rvsingle.dp.rf.rf\[20\]\[0\] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10985_ _05423_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__clkbuf_1
X_12724_ clknet_leaf_61_clk _00182_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12655_ clknet_leaf_36_clk _00113_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11606_ _05764_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12586_ clknet_leaf_83_clk _00044_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11537_ _05721_ _05722_ _05723_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold409 rvsingle.dp.rf.rf\[8\]\[24\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
X_11468_ _05685_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__clkbuf_1
X_13207_ clknet_leaf_64_clk _00665_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10419_ _04886_ net693 _05082_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11399_ _05322_ rvsingle.dp.rf.rf\[13\]\[2\] _05646_ VGND VGND VPWR VPWR _05648_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ clknet_leaf_40_clk _00596_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ clknet_leaf_43_clk _00527_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
X_07630_ _01419_ rvsingle.dp.rf.rf\[28\]\[4\] VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__or2_1
X_07561_ rvsingle.dp.rf.rf\[1\]\[4\] _02481_ _01496_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09300_ _04165_ _02101_ _04166_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__nand3_1
X_06512_ _01299_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__buf_8
X_07492_ _02408_ _02409_ _02410_ _02412_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09231_ _04148_ _04149_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__nand2_1
X_06443_ _01202_ _01364_ _01231_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06374_ _01295_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__clkbuf_8
X_09162_ _01225_ rvsingle.dp.rf.rf\[30\]\[31\] VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08113_ _01650_ rvsingle.dp.rf.rf\[26\]\[1\] _01104_ _03033_ VGND VGND VPWR VPWR
+ _03034_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_114_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09093_ _04008_ _04012_ _01189_ _02469_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__a31o_2
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08044_ _01067_ _01081_ _02914_ _02913_ _01083_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09995_ _04807_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__clkbuf_4
X_08946_ _01127_ rvsingle.dp.rf.rf\[10\]\[25\] VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__nor2_1
X_08877_ _01677_ rvsingle.dp.rf.rf\[3\]\[24\] _03797_ VGND VGND VPWR VPWR _03798_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07828_ _02375_ _02748_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07759_ _02677_ _02679_ _02291_ _01217_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__a31oi_1
X_10770_ _05292_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09429_ _04247_ _04332_ _04336_ _04337_ VGND VGND VPWR VPWR DataAdr[3] sky130_fd_sc_hd__o22ai_4
XFILLER_0_164_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12440_ clknet_leaf_34_clk _00924_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[27\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12371_ clknet_leaf_29_clk _00855_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11322_ net124 _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11253_ _05314_ _05566_ _05567_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__a21oi_1
X_10204_ _04738_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__buf_2
X_11184_ _05529_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10135_ _04738_ _04739_ _04927_ _04928_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__or4_4
X_10066_ _04425_ _04866_ _04867_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10968_ _05412_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12707_ clknet_leaf_124_clk _00165_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10899_ _05372_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__buf_6
XFILLER_0_54_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12638_ clknet_leaf_150_clk _00096_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ clknet_leaf_16_clk _01053_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold206 rvsingle.dp.rf.rf\[1\]\[22\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold217 rvsingle.dp.rf.rf\[19\]\[16\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 rvsingle.dp.rf.rf\[2\]\[28\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 rvsingle.dp.rf.rf\[4\]\[29\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ rvsingle.dp.rf.rf\[0\]\[15\] rvsingle.dp.rf.rf\[1\]\[15\] _02440_ VGND VGND
+ VPWR VPWR _03721_ sky130_fd_sc_hd__mux2_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ PC[23] _04612_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__xnor2_4
X_06992_ _01208_ _01908_ _01910_ _01912_ _01222_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__o221ai_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ rvsingle.dp.rf.rf\[19\]\[15\] _02478_ _01490_ VGND VGND VPWR VPWR _03652_
+ sky130_fd_sc_hd__o21ai_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08662_ _02929_ rvsingle.dp.rf.rf\[7\]\[14\] _01427_ _03582_ VGND VGND VPWR VPWR
+ _03583_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07613_ _02530_ _02533_ _01591_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__a21oi_2
X_08593_ _02117_ rvsingle.dp.rf.rf\[8\]\[12\] _01530_ VGND VGND VPWR VPWR _03514_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_72_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07544_ _01450_ _02293_ _01247_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07475_ _01847_ rvsingle.dp.rf.rf\[22\]\[6\] VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09214_ _04060_ _04062_ _01250_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__a21boi_2
X_06426_ _01288_ _01290_ _01347_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09145_ _01196_ rvsingle.dp.rf.rf\[12\]\[31\] VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06357_ _01139_ rvsingle.dp.rf.rf\[26\]\[29\] _01261_ VGND VGND VPWR VPWR _01280_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09076_ rvsingle.dp.rf.rf\[9\]\[26\] _01297_ _01310_ _03995_ VGND VGND VPWR VPWR
+ _03996_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_4_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06288_ _01204_ _01205_ _01210_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08027_ _02944_ _02945_ _01172_ _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__o211ai_1
Xhold740 rvsingle.dp.rf.rf\[29\]\[4\] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 rvsingle.dp.rf.rf\[4\]\[9\] VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold762 rvsingle.dp.rf.rf\[26\]\[1\] VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 rvsingle.dp.rf.rf\[21\]\[29\] VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold784 rvsingle.dp.rf.rf\[23\]\[27\] VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 rvsingle.dp.rf.rf\[16\]\[1\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ DataAdr[12] ReadData[12] _04750_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__mux2_1
X_08929_ rvsingle.dp.rf.rf\[19\]\[25\] _03839_ _03840_ VGND VGND VPWR VPWR _03850_
+ sky130_fd_sc_hd__o21ai_1
X_11940_ _05934_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ reset VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__buf_4
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10822_ _05085_ _05324_ _05325_ net118 VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10753_ _04782_ net583 _05274_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10684_ _04786_ rvsingle.dp.rf.rf\[21\]\[10\] _05235_ VGND VGND VPWR VPWR _05245_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12423_ clknet_leaf_99_clk _00907_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12354_ _05763_ net221 _06121_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__mux2_1
X_11305_ _05595_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12285_ _06091_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__clkbuf_1
X_11236_ _05557_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__clkbuf_1
X_11167_ _05307_ net451 _05511_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__mux2_1
X_10118_ _04909_ _04913_ _04729_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__o21ai_1
X_11098_ _05481_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__clkbuf_1
X_10049_ _04853_ net304 _04847_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07260_ _01450_ _02168_ _02180_ _01247_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__o211a_4
XFILLER_0_144_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06211_ Instr[20] VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_170_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07191_ _02108_ _02109_ _01503_ _02111_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06142_ _01065_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__buf_4
XFILLER_0_170_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09901_ _04727_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09832_ PC[25] PC[26] _04639_ PC[27] VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _04589_ _04592_ _04591_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__a21oi_1
X_06975_ _01875_ _01884_ _01682_ _01895_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__o211ai_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _01545_ rvsingle.dp.rf.rf\[2\]\[14\] _02337_ _03634_ VGND VGND VPWR VPWR
+ _03635_ sky130_fd_sc_hd__o211ai_1
X_09694_ _01225_ _04505_ _04506_ _04507_ PC[15] VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__a311o_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _01303_ _01351_ _03512_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__o21ai_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _03487_ _03489_ _01315_ _03496_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__o211a_2
XFILLER_0_77_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07527_ _01229_ _02441_ _02446_ _02447_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_147_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07458_ _01086_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06409_ _01330_ rvsingle.dp.rf.rf\[30\]\[29\] VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07389_ _02308_ _01730_ _01427_ _02309_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09128_ _01133_ _04042_ _04047_ _01117_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_33_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09059_ Instr[31] _01961_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12070_ _05137_ _05167_ _05976_ net358 VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__a2bb2o_1
Xhold570 rvsingle.dp.rf.rf\[2\]\[10\] VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 rvsingle.dp.rf.rf\[25\]\[0\] VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 rvsingle.dp.rf.rf\[9\]\[12\] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _05418_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__buf_8
X_12972_ clknet_leaf_52_clk _00430_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ _04852_ net230 _05924_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _05132_ net568 _05885_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__mux2_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _04909_ _04913_ _05271_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__o21ai_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11785_ _05132_ net352 _05845_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10736_ _05273_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__buf_8
XFILLER_0_103_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10667_ _05236_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12406_ clknet_leaf_31_clk _00890_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ clknet_leaf_82_clk _00814_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10598_ _05197_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12337_ _04839_ net700 _06110_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12268_ _06084_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__clkbuf_1
X_11219_ _05548_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12199_ _04904_ _04973_ _05316_ _06065_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__a31o_1
XFILLER_0_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06760_ _01670_ _01673_ _01634_ _01680_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_37_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06691_ _01611_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__clkbuf_8
X_08430_ _01768_ _03348_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nand3_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08361_ _03232_ _01537_ _03281_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07312_ _01512_ _02225_ _02227_ _01506_ _02232_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_128_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08292_ rvsingle.dp.rf.rf\[31\]\[10\] _01267_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__or2b_1
XFILLER_0_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07243_ _02163_ rvsingle.dp.rf.rf\[10\]\[17\] VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07174_ _02093_ _02094_ _01447_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09815_ _04644_ _04634_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__nor2_1
X_09746_ _04547_ _04560_ _04573_ _04578_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__or4_1
X_06958_ rvsingle.dp.rf.rf\[25\]\[22\] _01878_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ PC[12] _04500_ PC[13] VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__a21oi_1
X_06889_ rvsingle.dp.rf.rf\[11\]\[23\] _01441_ _01809_ VGND VGND VPWR VPWR _01810_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ rvsingle.dp.rf.rf\[29\]\[12\] _01492_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__or2b_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _01694_ _03474_ _03479_ _01699_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11570_ net160 _05726_ _05745_ _05737_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10521_ _04747_ rvsingle.dp.rf.rf\[9\]\[2\] _05152_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13240_ clknet_leaf_24_clk _00698_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10452_ _05111_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13171_ clknet_leaf_48_clk _00629_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10383_ _05073_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__clkbuf_1
X_12122_ _06009_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__buf_6
XFILLER_0_130_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12053_ _04833_ net470 _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11004_ _05209_ rvsingle.dp.rf.rf\[31\]\[13\] _05431_ VGND VGND VPWR VPWR _05434_
+ sky130_fd_sc_hd__mux2_1
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ clknet_leaf_141_clk _00413_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _04807_ net492 _05913_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__mux2_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 _06048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12886_ clknet_leaf_32_clk _00344_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _01148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_262 _01531_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11837_ _05344_ net333 _05874_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__mux2_1
XANTENNA_273 _01828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_284 _04817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 rvsingle.dp.rf.rf\[8\]\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11768_ _05846_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10719_ _05263_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11699_ _04801_ net493 _05806_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_991 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13369_ clknet_leaf_16_clk _00797_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07930_ _02848_ _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__nand2_4
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07861_ rvsingle.dp.rf.rf\[27\]\[2\] _01381_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__or2b_1
X_09600_ _04139_ _04363_ _04426_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__o21a_2
X_06812_ _01295_ rvsingle.dp.rf.rf\[31\]\[20\] _01732_ VGND VGND VPWR VPWR _01733_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07792_ _01125_ rvsingle.dp.rf.rf\[2\]\[3\] _01647_ _02712_ VGND VGND VPWR VPWR _02713_
+ sky130_fd_sc_hd__o211ai_1
X_09531_ _04219_ VGND VGND VPWR VPWR DataAdr[20] sky130_fd_sc_hd__inv_6
X_06743_ _01653_ _01663_ _01526_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__nand3_1
XFILLER_0_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09462_ _04140_ net825 _01067_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__o21ai_2
X_06674_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__buf_8
X_08413_ _01105_ _03330_ _03331_ _02483_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09393_ _04155_ _03054_ _04157_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08344_ _01558_ rvsingle.dp.rf.rf\[26\]\[8\] _01777_ VGND VGND VPWR VPWR _03265_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_171_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08275_ rvsingle.dp.rf.rf\[17\]\[10\] _01743_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07226_ _02143_ _02144_ _02146_ _01565_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_144_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07157_ rvsingle.dp.rf.rf\[12\]\[18\] rvsingle.dp.rf.rf\[13\]\[18\] _01432_ VGND
+ VGND VPWR VPWR _02078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07088_ _01634_ _02002_ _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__nand3_2
XFILLER_0_121_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09729_ _01224_ _02912_ _01175_ _04507_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__a31o_1
X_12740_ clknet_leaf_102_clk _00198_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ clknet_leaf_2_clk _00129_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11622_ _05724_ net563 _05775_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11553_ net113 _05731_ _05735_ _05157_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10504_ net77 VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11484_ _05693_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13223_ clknet_leaf_101_clk _00681_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10435_ _04724_ _04927_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13154_ clknet_leaf_128_clk _00612_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10366_ _04965_ _04927_ _05063_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__or3_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _06022_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__clkbuf_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13085_ clknet_leaf_146_clk _00543_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _04755_ net786 _05022_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__mux2_1
X_12036_ _05986_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ clknet_leaf_81_clk _00396_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ clknet_leaf_114_clk _00327_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06390_ _01195_ rvsingle.dp.rf.rf\[0\]\[29\] VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08060_ _01229_ _02975_ _02980_ _02447_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07011_ rvsingle.dp.rf.rf\[20\]\[19\] rvsingle.dp.rf.rf\[21\]\[19\] rvsingle.dp.rf.rf\[22\]\[19\]
+ rvsingle.dp.rf.rf\[23\]\[19\] _01463_ _01456_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08962_ rvsingle.dp.rf.rf\[20\]\[25\] rvsingle.dp.rf.rf\[21\]\[25\] rvsingle.dp.rf.rf\[22\]\[25\]
+ rvsingle.dp.rf.rf\[23\]\[25\] _01194_ _01201_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__mux4_1
X_07913_ _01462_ rvsingle.dp.rf.rf\[16\]\[2\] _01299_ VGND VGND VPWR VPWR _02834_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08893_ _01219_ _03809_ _01316_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07844_ _02763_ _02764_ _02329_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07775_ _01188_ _02682_ _02695_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09514_ _04377_ _02774_ _02797_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__and3_4
XFILLER_0_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06726_ _01103_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__buf_6
XFILLER_0_94_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09445_ _02534_ _02573_ _04350_ _04347_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__o211ai_2
X_06657_ _01536_ _01537_ _01153_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__nand4_2
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09376_ _01837_ _01581_ _02067_ _04123_ _04291_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a311o_1
XFILLER_0_163_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06588_ _01508_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08327_ _03244_ _03245_ _03247_ _02483_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_164_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08258_ _01136_ rvsingle.dp.rf.rf\[12\]\[10\] _01519_ VGND VGND VPWR VPWR _03179_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07209_ rvsingle.dp.rf.rf\[11\]\[17\] _02030_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08189_ _03092_ _03098_ _01377_ _03109_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10220_ _04980_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__clkbuf_1
X_10151_ _04778_ rvsingle.dp.rf.rf\[28\]\[8\] _04930_ VGND VGND VPWR VPWR _04938_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10082_ _04879_ _04880_ _04881_ ReadData[27] _04715_ VGND VGND VPWR VPWR _04882_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10984_ _05377_ rvsingle.dp.rf.rf\[31\]\[4\] _05419_ VGND VGND VPWR VPWR _05423_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12723_ clknet_leaf_27_clk _00181_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12654_ clknet_leaf_72_clk _00112_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11605_ _05763_ net442 _05729_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12585_ clknet_leaf_97_clk _00043_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11536_ _04976_ _05417_ _05149_ _02873_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__o31a_1
XFILLER_0_81_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11467_ _05318_ net681 _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13206_ clknet_leaf_64_clk _00664_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10418_ _05090_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11398_ _05647_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__clkbuf_1
X_13137_ clknet_leaf_48_clk _00595_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _04892_ net297 _05044_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ clknet_leaf_51_clk _00526_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _05728_ net607 _05976_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__mux2_1
X_07560_ _01645_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06511_ _01426_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07491_ rvsingle.dp.rf.rf\[15\]\[6\] _01508_ _02411_ VGND VGND VPWR VPWR _02412_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09230_ _03573_ _03735_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__nor2_1
X_06442_ rvsingle.dp.rf.rf\[2\]\[28\] rvsingle.dp.rf.rf\[3\]\[28\] _01338_ VGND VGND
+ VPWR VPWR _01364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09161_ rvsingle.dp.rf.rf\[29\]\[31\] _01298_ _01311_ _04080_ VGND VGND VPWR VPWR
+ _04081_ sky130_fd_sc_hd__o211a_1
X_06373_ _01294_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__buf_6
XFILLER_0_145_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08112_ rvsingle.dp.rf.rf\[27\]\[1\] _01124_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09092_ _01231_ _04009_ _04011_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08043_ _02885_ _01481_ _01592_ _02906_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__nand4_2
XFILLER_0_114_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09994_ _04365_ _04805_ _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_0_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08945_ _03863_ _03782_ _03865_ _01506_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__a31o_1
X_08876_ _01255_ rvsingle.dp.rf.rf\[2\]\[24\] _01530_ VGND VGND VPWR VPWR _03797_
+ sky130_fd_sc_hd__o21a_1
X_07827_ Instr[10] _01078_ _02697_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__o21a_2
XFILLER_0_98_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07758_ _02271_ rvsingle.dp.rf.rf\[15\]\[3\] _01300_ _02678_ VGND VGND VPWR VPWR
+ _02679_ sky130_fd_sc_hd__o211ai_1
X_06709_ _01557_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07689_ _01862_ rvsingle.dp.rf.rf\[10\]\[5\] VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09428_ _02751_ _02856_ _04335_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09359_ _02100_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12370_ clknet_leaf_57_clk _00854_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11321_ _04916_ _04918_ _04728_ _04922_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__and4b_2
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11252_ net142 _05566_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10203_ _04965_ _04927_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__nor2_1
X_11183_ _05318_ net766 _05528_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10134_ _04713_ _04724_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__nand2_4
X_10065_ _04425_ _04643_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10967_ _05187_ net385 _05401_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ clknet_leaf_131_clk _00164_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10898_ _04738_ _04733_ _05371_ _04739_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__or4b_4
XFILLER_0_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12637_ clknet_leaf_144_clk _00095_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12568_ clknet_leaf_22_clk _01052_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11519_ _05407_ net556 _05706_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12499_ clknet_leaf_33_clk _00983_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold207 rvsingle.dp.rf.rf\[3\]\[22\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 rvsingle.dp.rf.rf\[8\]\[11\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 rvsingle.dp.rf.rf\[26\]\[24\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _01911_ _01309_ _01711_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__a21o_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _01595_ rvsingle.dp.rf.rf\[18\]\[15\] VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__nor2_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _01425_ rvsingle.dp.rf.rf\[6\]\[14\] VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__or2_1
X_07612_ _01178_ _02532_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__nand2_1
X_08592_ _01452_ _03497_ _03512_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07543_ _02430_ _02432_ _02463_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__nand3_4
XFILLER_0_72_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07474_ _01091_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09213_ _04131_ _01066_ _04123_ _04113_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__a211o_2
X_06425_ _01248_ _01324_ _01346_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__and3_2
XFILLER_0_147_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09144_ rvsingle.dp.rf.rf\[8\]\[31\] rvsingle.dp.rf.rf\[9\]\[31\] rvsingle.dp.rf.rf\[10\]\[31\]
+ rvsingle.dp.rf.rf\[11\]\[31\] _01196_ _01203_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__mux4_1
X_06356_ _01276_ _01094_ _01134_ _01278_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_44_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09075_ _01330_ rvsingle.dp.rf.rf\[8\]\[26\] VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__or2_1
X_06287_ _01209_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_170_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08026_ rvsingle.dp.rf.rf\[13\]\[0\] _01423_ _01307_ _02946_ VGND VGND VPWR VPWR
+ _02947_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold730 rvsingle.dp.rf.rf\[27\]\[15\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 rvsingle.dp.rf.rf\[15\]\[5\] VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold752 rvsingle.dp.rf.rf\[29\]\[5\] VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 rvsingle.dp.rf.rf\[27\]\[13\] VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 rvsingle.dp.rf.rf\[28\]\[4\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 rvsingle.dp.rf.rf\[14\]\[17\] VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 rvsingle.dp.rf.rf\[29\]\[11\] VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd3_1
X_09977_ _04792_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08928_ _01257_ rvsingle.dp.rf.rf\[18\]\[25\] VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__nor2_1
X_08859_ rvsingle.dp.rf.rf\[23\]\[24\] _03778_ _03779_ VGND VGND VPWR VPWR _03780_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _05896_ _05860_ _05897_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10821_ _05320_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__clkbuf_8
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10752_ _05282_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10683_ _05244_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12422_ clknet_leaf_108_clk _00906_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12353_ _06128_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11304_ _05354_ rvsingle.dp.rf.rf\[15\]\[24\] _05591_ VGND VGND VPWR VPWR _05595_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12284_ _05763_ net264 _06073_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__mux2_1
X_11235_ _05304_ net800 _05552_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__mux2_1
X_11166_ _05518_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__clkbuf_1
X_10117_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__clkbuf_4
X_11097_ _05307_ net606 _05469_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__mux2_1
X_10048_ _04852_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_171_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold90 rvsingle.dp.rf.rf\[5\]\[31\] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11999_ _05966_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06210_ _01133_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07190_ rvsingle.dp.rf.rf\[31\]\[17\] _01861_ _02110_ VGND VGND VPWR VPWR _02111_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06141_ _01064_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09900_ Instr[7] Instr[8] VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__and2b_1
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09831_ PC[25] PC[26] PC[27] _04639_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__and4_2
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06974_ _01157_ _01889_ _01894_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__nand3_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ Instr[31] PC[21] VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__xnor2_2
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ rvsingle.dp.rf.rf\[3\]\[14\] _01877_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__or2b_1
X_09693_ _04536_ PC[15] VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08644_ _03513_ _03562_ _03564_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__nand3_4
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _01422_ _03490_ _03495_ _01221_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_77_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07526_ _01216_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__buf_6
XFILLER_0_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07457_ _01763_ rvsingle.dp.rf.rf\[26\]\[6\] VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06408_ _01329_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07388_ _01468_ rvsingle.dp.rf.rf\[20\]\[7\] VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09127_ _01106_ _04044_ _04046_ _01132_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_33_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06339_ rvsingle.dp.rf.rf\[4\]\[29\] rvsingle.dp.rf.rf\[5\]\[29\] rvsingle.dp.rf.rf\[6\]\[29\]
+ rvsingle.dp.rf.rf\[7\]\[29\] _01257_ _01261_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__mux4_1
X_09058_ _01153_ _03956_ _03977_ _01482_ _01184_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__a41o_1
X_08009_ _01240_ rvsingle.dp.rf.rf\[18\]\[0\] _01197_ VGND VGND VPWR VPWR _02930_
+ sky130_fd_sc_hd__o21a_1
Xhold560 rvsingle.dp.rf.rf\[4\]\[10\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold571 rvsingle.dp.rf.rf\[20\]\[21\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ _05442_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__clkbuf_1
Xhold582 rvsingle.dp.rf.rf\[2\]\[23\] VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 rvsingle.dp.rf.rf\[30\]\[13\] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ clknet_leaf_86_clk _00429_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _05925_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__clkbuf_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _05888_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ net47 VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__inv_2
X_11784_ _05851_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__clkbuf_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_898 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10735_ _04917_ _04920_ _04921_ _04915_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10666_ _04736_ net499 _05235_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12405_ clknet_leaf_36_clk _00889_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_13385_ clknet_leaf_94_clk _00813_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10597_ _04755_ net802 _05194_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12336_ _06119_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12267_ _05173_ net494 _06073_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11218_ _05476_ net668 _05541_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__mux2_1
X_12198_ _04982_ _04983_ _04981_ _05003_ net313 VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__o41a_1
X_11149_ _05439_ rvsingle.dp.rf.rf\[16\]\[18\] _05499_ VGND VGND VPWR VPWR _05510_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06690_ _01610_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08360_ _03255_ _01083_ _02505_ _03280_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__nand4_4
XFILLER_0_86_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07311_ _02228_ _02229_ _01112_ _02231_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_86_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08291_ rvsingle.dp.rf.rf\[29\]\[10\] _02005_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07242_ _01190_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__buf_4
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07173_ rvsingle.dp.rf.rf\[28\]\[18\] rvsingle.dp.rf.rf\[29\]\[18\] rvsingle.dp.rf.rf\[30\]\[18\]
+ rvsingle.dp.rf.rf\[31\]\[18\] _01241_ _01199_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09814_ _04398_ _04643_ _04647_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[25\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09745_ _04398_ _04580_ _04584_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[19\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06957_ _01877_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _01726_ rvsingle.dp.rf.rf\[10\]\[23\] _01808_ VGND VGND VPWR VPWR _01809_
+ sky130_fd_sc_hd__o21a_1
X_09676_ _04521_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__clkbuf_2
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _03539_ _03542_ _01156_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__o211ai_2
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08558_ _03475_ _03476_ _03477_ _03478_ _01702_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_154_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07509_ _02428_ _01183_ _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__nand3_1
XFILLER_0_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08489_ rvsingle.dp.rf.rf\[25\]\[13\] _01136_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10520_ _05153_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_959 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10451_ _04774_ rvsingle.dp.rf.rf\[24\]\[7\] _05110_ VGND VGND VPWR VPWR _05111_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13170_ clknet_leaf_51_clk _00628_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10382_ _04778_ rvsingle.dp.rf.rf\[25\]\[8\] _05071_ VGND VGND VPWR VPWR _05073_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12121_ _06030_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12052_ _05975_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__buf_6
Xhold390 rvsingle.dp.rf.rf\[8\]\[6\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _05433_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__clkbuf_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ clknet_leaf_1_clk _00412_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _05916_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__clkbuf_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _05469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12885_ clknet_leaf_36_clk _00343_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_241 _06048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_252 _01255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 _01539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11836_ _05879_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _01853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 _04817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_296 rvsingle.dp.rf.rf\[8\]\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11767_ _04795_ net251 _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__mux2_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10718_ _04877_ net756 _05257_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11698_ _05808_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10649_ _05225_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13368_ clknet_leaf_20_clk _00796_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12319_ _05744_ net284 _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13299_ clknet_leaf_68_clk _00757_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07860_ rvsingle.dp.rf.rf\[25\]\[2\] _01613_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__and2b_1
X_06811_ _01462_ rvsingle.dp.rf.rf\[30\]\[20\] _01198_ VGND VGND VPWR VPWR _01732_
+ sky130_fd_sc_hd__o21a_1
X_07791_ rvsingle.dp.rf.rf\[3\]\[3\] _01606_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__or2b_1
XFILLER_0_64_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06742_ _01655_ _01657_ _01659_ _01600_ _01662_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__o311ai_1
X_09530_ _04284_ VGND VGND VPWR VPWR DataAdr[19] sky130_fd_sc_hd__inv_2
XFILLER_0_78_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09461_ _02914_ _02913_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__nand2_1
X_06673_ _01095_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__buf_6
X_08412_ _01513_ rvsingle.dp.rf.rf\[2\]\[9\] _02059_ _03332_ VGND VGND VPWR VPWR _03333_
+ sky130_fd_sc_hd__o211ai_1
X_09392_ _04301_ _04302_ _04305_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__and4_1
X_08343_ _03262_ _01744_ _03263_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08274_ _01268_ rvsingle.dp.rf.rf\[16\]\[10\] VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07225_ rvsingle.dp.rf.rf\[1\]\[17\] _01842_ _01092_ _02145_ VGND VGND VPWR VPWR
+ _02146_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_117_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07156_ _01943_ rvsingle.dp.rf.rf\[15\]\[18\] _01451_ _02076_ VGND VGND VPWR VPWR
+ _02077_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07087_ _01092_ _02003_ _02004_ _01617_ _02007_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07989_ Instr[2] VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__clkbuf_4
X_09728_ _04561_ _04559_ _04568_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09659_ _01175_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__clkbuf_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ clknet_leaf_150_clk _00128_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _05774_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11552_ _04759_ _05732_ _05733_ _05060_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__and4_1
XFILLER_0_65_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10503_ _05139_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11483_ _05428_ net467 _05684_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13222_ clknet_leaf_91_clk _00680_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_10434_ _04719_ _05098_ _05100_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13153_ clknet_leaf_140_clk _00611_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10365_ Instr[8] _04732_ Instr[7] VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__or3b_1
XFILLER_0_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _05744_ net450 _06019_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__mux2_1
X_13084_ clknet_leaf_151_clk _00542_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10296_ _05024_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__clkbuf_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12035_ _04785_ net613 _05983_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12937_ clknet_leaf_97_clk _00395_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ clknet_leaf_107_clk _00326_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11819_ _05870_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__clkbuf_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12799_ clknet_leaf_1_clk _00257_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07010_ _01590_ _01742_ _01840_ _01930_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__nor4_2
XFILLER_0_3_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08961_ _01837_ _01581_ _03879_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07912_ _01420_ rvsingle.dp.rf.rf\[18\]\[2\] _01696_ _02832_ VGND VGND VPWR VPWR
+ _02833_ sky130_fd_sc_hd__o211ai_1
X_08892_ _01722_ _03810_ _01478_ _03812_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07843_ rvsingle.dp.rf.rf\[1\]\[2\] _01613_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__and2b_1
X_07774_ _02686_ _02688_ _01187_ _02694_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__o211ai_4
X_09513_ _04392_ VGND VGND VPWR VPWR WriteData[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06725_ _01645_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06656_ _01378_ _01556_ _01576_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__nand3_2
X_09444_ _03056_ _04347_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__a21o_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09375_ _02081_ _02097_ _02068_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__o21a_1
X_06587_ _01086_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08326_ rvsingle.dp.rf.rf\[1\]\[8\] _02478_ _02395_ _03246_ VGND VGND VPWR VPWR _03247_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08257_ rvsingle.dp.rf.rf\[15\]\[10\] _01769_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_668 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07208_ _01126_ rvsingle.dp.rf.rf\[10\]\[17\] VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08188_ _03103_ _03108_ _01505_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__nand3_2
X_07139_ _01268_ rvsingle.dp.rf.rf\[10\]\[18\] _02059_ VGND VGND VPWR VPWR _02060_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10150_ _04937_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10081_ _02910_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_148_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_148_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10983_ _05422_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12722_ clknet_leaf_47_clk _00180_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12653_ clknet_leaf_43_clk _00111_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11604_ _04891_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__buf_2
XFILLER_0_81_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12584_ clknet_leaf_123_clk _00042_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11535_ _04720_ _05142_ _04967_ _04968_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__and4_1
XFILLER_0_151_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11466_ _05683_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__buf_6
XFILLER_0_123_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13205_ clknet_leaf_24_clk _00663_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10417_ _04877_ net769 _05082_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11397_ _05318_ rvsingle.dp.rf.rf\[13\]\[1\] _05646_ VGND VGND VPWR VPWR _05647_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13136_ clknet_leaf_71_clk _00594_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _05051_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _04892_ net289 _05001_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__mux2_1
X_13067_ clknet_leaf_90_clk _00525_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12018_ _05977_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_139_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_139_clk sky130_fd_sc_hd__clkbuf_16
X_06510_ _01230_ _01418_ _01430_ _01222_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__o211ai_1
X_07490_ _01267_ rvsingle.dp.rf.rf\[14\]\[6\] _01489_ VGND VGND VPWR VPWR _02411_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06441_ rvsingle.dp.rf.rf\[1\]\[28\] _01298_ _01311_ _01362_ VGND VGND VPWR VPWR
+ _01363_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_111_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09160_ _01225_ rvsingle.dp.rf.rf\[28\]\[31\] VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06372_ _01293_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08111_ rvsingle.dp.rf.rf\[25\]\[1\] _01381_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09091_ _02191_ _04010_ _01218_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08042_ _01870_ _02915_ _02962_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09993_ _01169_ _02259_ _01170_ _04534_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__or4b_2
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08944_ _03778_ rvsingle.dp.rf.rf\[5\]\[25\] _03864_ VGND VGND VPWR VPWR _03865_
+ sky130_fd_sc_hd__o21ai_1
X_08875_ rvsingle.dp.rf.rf\[0\]\[24\] rvsingle.dp.rf.rf\[1\]\[24\] _02117_ VGND VGND
+ VPWR VPWR _03796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07826_ _01065_ _01074_ _01481_ _02698_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__o221a_1
XFILLER_0_169_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07757_ _01419_ rvsingle.dp.rf.rf\[14\]\[3\] VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06708_ _01518_ rvsingle.dp.rf.rf\[6\]\[20\] _01620_ VGND VGND VPWR VPWR _01629_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07688_ _02375_ Instr[25] VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__nand2_2
X_09427_ _04333_ _04335_ _04135_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06639_ _01559_ rvsingle.dp.rf.rf\[0\]\[21\] VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09358_ _04249_ _04256_ _04268_ _04273_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__nand4_1
XFILLER_0_35_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08309_ _02469_ _03228_ _03229_ _03143_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_118_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09289_ _01585_ _01180_ _01586_ _01582_ _04143_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11320_ _05602_ _05566_ _05603_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11251_ _05417_ _05565_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__nor2_2
XFILLER_0_105_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10202_ _04724_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__clkbuf_4
X_11182_ _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__buf_6
X_10133_ _04722_ _04723_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__nand2_4
XFILLER_0_100_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10064_ _02908_ DataAdr[25] _04865_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10966_ _05411_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12705_ clknet_leaf_125_clk _00163_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10897_ _05370_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12636_ clknet_leaf_151_clk _00094_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12567_ clknet_leaf_16_clk _01051_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11518_ _05711_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12498_ clknet_leaf_36_clk _00982_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold208 rvsingle.dp.rf.rf\[17\]\[21\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold219 rvsingle.dp.rf.rf\[0\]\[29\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11449_ _05407_ net645 _05668_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ clknet_leaf_133_clk _00577_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ rvsingle.dp.rf.rf\[24\]\[22\] rvsingle.dp.rf.rf\[25\]\[22\] _01695_ VGND
+ VGND VPWR VPWR _01911_ sky130_fd_sc_hd__mux2_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ rvsingle.dp.rf.rf\[4\]\[14\] rvsingle.dp.rf.rf\[5\]\[14\] _01468_ VGND VGND
+ VPWR VPWR _03581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07611_ Instr[11] _01078_ _02531_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__o21a_1
X_08591_ _03501_ _03503_ _02315_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07542_ _02315_ _02449_ _02462_ _01246_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07473_ _01490_ _02390_ _02391_ _01564_ _02393_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_64_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09212_ _04110_ _04112_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__nand2_1
X_06424_ _01317_ _01334_ _01345_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__or3_1
XFILLER_0_146_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06355_ _01089_ rvsingle.dp.rf.rf\[23\]\[29\] _01107_ _01277_ VGND VGND VPWR VPWR
+ _01278_ sky130_fd_sc_hd__o211a_1
X_09143_ _04060_ _04062_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__nand2_4
XFILLER_0_115_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09074_ _01194_ rvsingle.dp.rf.rf\[10\]\[26\] _03993_ VGND VGND VPWR VPWR _03994_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06286_ _01208_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08025_ _01327_ rvsingle.dp.rf.rf\[12\]\[0\] VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold720 rvsingle.dp.rf.rf\[13\]\[15\] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 rvsingle.dp.rf.rf\[24\]\[3\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold742 rvsingle.dp.rf.rf\[28\]\[24\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold753 rvsingle.dp.rf.rf\[13\]\[7\] VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 rvsingle.dp.rf.rf\[25\]\[12\] VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 rvsingle.dp.rf.rf\[3\]\[2\] VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 rvsingle.dp.rf.rf\[26\]\[3\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 rvsingle.dp.rf.rf\[27\]\[8\] VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ _04790_ net339 _04791_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__mux2_1
X_08927_ _01106_ _03844_ _03845_ _03846_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_157_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08858_ _01643_ rvsingle.dp.rf.rf\[22\]\[24\] _01648_ VGND VGND VPWR VPWR _03779_
+ sky130_fd_sc_hd__o21a_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07809_ _01797_ rvsingle.dp.rf.rf\[26\]\[3\] _01647_ _02729_ VGND VGND VPWR VPWR
+ _02730_ sky130_fd_sc_hd__o211ai_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ rvsingle.dp.rf.rf\[19\]\[15\] _01424_ _03709_ VGND VGND VPWR VPWR _03710_
+ sky130_fd_sc_hd__o21ai_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10820_ _04982_ _04983_ _04981_ _04754_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__or4b_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10751_ _04778_ rvsingle.dp.rf.rf\[20\]\[8\] _05274_ VGND VGND VPWR VPWR _05282_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10682_ _04782_ net325 _05235_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12421_ clknet_leaf_114_clk _00905_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12352_ _04885_ net305 _06121_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11303_ _05594_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__clkbuf_1
X_12283_ _04886_ _05183_ _05832_ _06090_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11234_ _05556_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__clkbuf_1
X_11165_ _05407_ rvsingle.dp.rf.rf\[16\]\[26\] _05511_ VGND VGND VPWR VPWR _05518_
+ sky130_fd_sc_hd__mux2_1
X_10116_ _01169_ _02259_ _01170_ _04910_ _04911_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__o32a_2
X_11096_ _05460_ net179 _05182_ _05464_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10047_ _04365_ _04850_ _04851_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__o21ai_4
Xhold80 rvsingle.dp.rf.rf\[29\]\[31\] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 rvsingle.dp.rf.rf\[7\]\[9\] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11998_ _04869_ net293 _05960_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10949_ _05402_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12619_ clknet_leaf_64_clk _00077_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06140_ Instr[30] Instr[5] _01059_ _01060_ _01063_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09830_ _04367_ _04654_ _04660_ _04662_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[26\]
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _04597_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__or2_2
X_06973_ _01890_ _01891_ _01503_ _01893_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__o211ai_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ rvsingle.dp.rf.rf\[1\]\[14\] _03258_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__and2b_1
X_09692_ _01225_ _04505_ _04506_ _04507_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__a31o_1
X_08643_ _02473_ _02102_ _03142_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08574_ _03491_ _03492_ _02543_ _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__o211ai_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07525_ _02442_ _02443_ _02444_ _02445_ _02273_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07456_ _02376_ _02372_ _01485_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06407_ _01328_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__buf_8
XFILLER_0_91_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07387_ rvsingle.dp.rf.rf\[21\]\[7\] VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09126_ _01488_ rvsingle.dp.rf.rf\[27\]\[26\] _01491_ _04045_ VGND VGND VPWR VPWR
+ _04046_ sky130_fd_sc_hd__o211ai_1
X_06338_ _01260_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09057_ _03961_ _03966_ _03976_ _01378_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__o211ai_4
X_06269_ _01191_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08008_ _01293_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__clkbuf_8
Xhold550 rvsingle.dp.rf.rf\[10\]\[26\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold561 rvsingle.dp.rf.rf\[6\]\[15\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 rvsingle.dp.rf.rf\[16\]\[2\] VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 rvsingle.dp.rf.rf\[20\]\[9\] VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold594 rvsingle.dp.rf.rf\[18\]\[27\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ _04777_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__clkbuf_4
X_12970_ clknet_leaf_81_clk _00428_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _04845_ net384 _05924_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11852_ _05757_ net256 _05885_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__mux2_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _05311_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__clkbuf_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _05757_ rvsingle.dp.rf.rf\[7\]\[23\] _05845_ VGND VGND VPWR VPWR _05851_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10734_ _04719_ _05271_ _05272_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10665_ _05234_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__buf_8
X_12404_ clknet_leaf_21_clk _00888_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_13384_ clknet_leaf_122_clk _00812_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10596_ _05196_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12335_ _04833_ net651 _06110_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12266_ _06083_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11217_ _05547_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__clkbuf_1
X_12197_ _06064_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11148_ _05509_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__clkbuf_1
X_11079_ _05471_ _05474_ _05463_ net183 VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_37_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07310_ rvsingle.dp.rf.rf\[31\]\[16\] _01509_ _02230_ VGND VGND VPWR VPWR _02231_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08290_ _01878_ rvsingle.dp.rf.rf\[28\]\[10\] VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07241_ _01299_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07172_ _01460_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__buf_6
XFILLER_0_54_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09813_ _04366_ _04645_ _04646_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09744_ _04422_ _04423_ _04583_ _04427_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__o211a_1
X_06956_ _01095_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09675_ PC[12] PC[13] _04500_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__and3_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06887_ _01198_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__buf_6
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _01660_ _03543_ _03544_ _02351_ _03546_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__o311ai_2
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ rvsingle.dp.rf.rf\[5\]\[13\] _01901_ _02285_ VGND VGND VPWR VPWR _03478_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07508_ Instr[26] _01083_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08488_ _01607_ rvsingle.dp.rf.rf\[24\]\[13\] _01489_ VGND VGND VPWR VPWR _03409_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07439_ _02308_ _01614_ _02320_ _02359_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10450_ _05102_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__buf_8
XFILLER_0_135_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09109_ _04025_ _04026_ _02236_ _04028_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_21_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10381_ _05072_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__clkbuf_1
X_12120_ _04833_ net472 _06019_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12051_ _05993_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold380 rvsingle.dp.rf.rf\[13\]\[30\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 rvsingle.dp.rf.rf\[2\]\[27\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11002_ _05207_ rvsingle.dp.rf.rf\[31\]\[12\] _05431_ VGND VGND VPWR VPWR _05433_
+ sky130_fd_sc_hd__mux2_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ clknet_leaf_9_clk _00411_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _04801_ net703 _05913_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__mux2_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ clknet_leaf_25_clk _00342_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_220 _05085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_231 _05499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 _06049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11835_ _04813_ net675 _05874_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__mux2_1
XANTENNA_253 _01255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 _01660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_275 _01862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _04817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_297 _01247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11766_ _05836_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__buf_6
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10717_ _05262_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11697_ _04795_ net363 _05806_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10648_ _04877_ net546 _05219_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13367_ clknet_leaf_16_clk _00795_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10579_ _05185_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__clkbuf_1
X_12318_ _06098_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__buf_6
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13298_ clknet_leaf_67_clk _00756_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_950 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12249_ _06078_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06810_ rvsingle.dp.rf.rf\[28\]\[20\] rvsingle.dp.rf.rf\[29\]\[20\] _01730_ VGND
+ VGND VPWR VPWR _01731_ sky130_fd_sc_hd__mux2_1
X_07790_ rvsingle.dp.rf.rf\[1\]\[3\] _01566_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06741_ _01656_ rvsingle.dp.rf.rf\[26\]\[20\] _01660_ _01661_ VGND VGND VPWR VPWR
+ _01662_ sky130_fd_sc_hd__o211ai_1
X_09460_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__buf_4
X_06672_ _01376_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__buf_12
X_08411_ rvsingle.dp.rf.rf\[3\]\[9\] _01492_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__or2b_1
X_09391_ _03825_ _03803_ _04143_ _03826_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08342_ _01763_ rvsingle.dp.rf.rf\[24\]\[8\] _01604_ VGND VGND VPWR VPWR _03263_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_80_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08273_ _01593_ _03182_ _03193_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__nand3_2
XFILLER_0_74_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07224_ _01607_ rvsingle.dp.rf.rf\[0\]\[17\] VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07155_ _01336_ rvsingle.dp.rf.rf\[14\]\[18\] VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07086_ _01796_ rvsingle.dp.rf.rf\[5\]\[19\] _02006_ VGND VGND VPWR VPWR _02007_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07988_ Instr[3] VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__clkbuf_4
X_09727_ _04559_ PC[16] _04546_ _04558_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__a31o_1
X_06939_ _01086_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__clkbuf_8
X_09658_ _02912_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__buf_4
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08609_ _03528_ _03529_ _02410_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09589_ Instr[25] _04429_ _04439_ _04419_ _04438_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__o221a_1
XFILLER_0_139_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _04976_ _05417_ _05371_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__or3_2
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11551_ net86 _05731_ _05734_ _05157_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10502_ _04904_ net323 _05126_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11482_ _05692_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13221_ clknet_leaf_123_clk _00679_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10433_ _04970_ _05099_ net17 VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13152_ clknet_leaf_118_clk _00610_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10364_ _04719_ _05059_ _05062_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_131_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12103_ _06021_ _05060_ _04924_ _06010_ net15 VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__a32o_1
X_13083_ clknet_leaf_135_clk _00541_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10295_ _04747_ rvsingle.dp.rf.rf\[26\]\[2\] _05022_ VGND VGND VPWR VPWR _05024_
+ sky130_fd_sc_hd__mux2_1
X_12034_ _05976_ net152 _05116_ _05146_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ clknet_leaf_105_clk _00394_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ clknet_leaf_116_clk _00325_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _05381_ net778 _05863_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12798_ clknet_leaf_134_clk _00256_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11749_ _05838_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08960_ _01581_ _03879_ _01837_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
X_07911_ rvsingle.dp.rf.rf\[19\]\[2\] _01191_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__or2b_1
X_08891_ _01229_ _03811_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__or2_1
X_07842_ _01607_ rvsingle.dp.rf.rf\[0\]\[2\] _01489_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07773_ _02302_ _02689_ _02693_ _02438_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__o211ai_2
X_09512_ _04377_ _02721_ _02745_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__and3_4
X_06724_ _01086_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09443_ _02661_ _02667_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__nand2_1
X_06655_ _01157_ _01570_ _01575_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__nand3_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09374_ _04214_ _03765_ _04276_ _04125_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__a31o_1
X_06586_ _01269_ rvsingle.dp.rf.rf\[30\]\[21\] VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08325_ _02627_ rvsingle.dp.rf.rf\[0\]\[8\] VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08256_ _01780_ rvsingle.dp.rf.rf\[14\]\[10\] VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07207_ rvsingle.dp.rf.rf\[9\]\[17\] _01088_ _01668_ _02127_ VGND VGND VPWR VPWR
+ _02128_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08187_ _03104_ _03105_ _02329_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__o211ai_1
X_07138_ _01519_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07069_ _01655_ _01986_ _01987_ _01768_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10080_ _02799_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__buf_4
X_10982_ _04755_ rvsingle.dp.rf.rf\[31\]\[3\] _05419_ VGND VGND VPWR VPWR _05422_
+ sky130_fd_sc_hd__mux2_1
X_12721_ clknet_leaf_49_clk _00179_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12652_ clknet_leaf_49_clk _00110_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11603_ _05762_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12583_ clknet_leaf_101_clk _00041_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11534_ _04718_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11465_ _04738_ _04739_ _05565_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__or3_2
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13204_ clknet_leaf_55_clk _00662_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10416_ _05089_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11396_ _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__buf_6
XFILLER_0_150_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13135_ clknet_leaf_37_clk _00593_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10347_ _04886_ net382 _05044_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ clknet_leaf_82_clk _00524_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10278_ _05013_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__clkbuf_1
X_12017_ _05724_ net578 _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12919_ clknet_leaf_7_clk _00377_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06440_ _01195_ rvsingle.dp.rf.rf\[0\]\[28\] VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06371_ Instr[15] VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08110_ _01602_ rvsingle.dp.rf.rf\[24\]\[1\] VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09090_ rvsingle.dp.rf.rf\[20\]\[26\] rvsingle.dp.rf.rf\[21\]\[26\] rvsingle.dp.rf.rf\[22\]\[26\]
+ rvsingle.dp.rf.rf\[23\]\[26\] _01242_ _01200_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08041_ _01337_ _01451_ _01245_ _02939_ _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__o311a_1
XFILLER_0_141_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09992_ _02908_ DataAdr[14] _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08943_ _01098_ rvsingle.dp.rf.rf\[4\]\[25\] _01105_ VGND VGND VPWR VPWR _03864_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
X_08874_ rvsingle.dp.rf.rf\[4\]\[24\] rvsingle.dp.rf.rf\[5\]\[24\] rvsingle.dp.rf.rf\[6\]\[24\]
+ rvsingle.dp.rf.rf\[7\]\[24\] _01562_ _01655_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07825_ _02721_ _01082_ _01152_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__nand4_4
XFILLER_0_79_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07756_ rvsingle.dp.rf.rf\[13\]\[3\] _02288_ _01436_ _02676_ VGND VGND VPWR VPWR
+ _02677_ sky130_fd_sc_hd__o211ai_1
X_06707_ _01625_ _01098_ _01626_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_94_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07687_ _01450_ _02593_ _02607_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09426_ _02803_ _02851_ _04334_ _04151_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__o22ai_1
X_06638_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__buf_4
XFILLER_0_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09357_ _04269_ _04270_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__o21a_2
XFILLER_0_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06569_ _01489_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08308_ _01065_ _01074_ _01961_ _03111_ _01580_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__o221a_1
X_09288_ _01742_ _04167_ _01590_ _01739_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_74_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08239_ _03157_ _02291_ _03159_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__nand3_2
XFILLER_0_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11250_ _04928_ _04722_ _04723_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__or3b_4
XFILLER_0_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10201_ _04963_ _04923_ _04964_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11181_ _04919_ _04927_ _04928_ _04738_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__or4b_4
X_10132_ _04719_ _04923_ _04926_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10063_ _02909_ _02799_ _02910_ ReadData[25] _04245_ VGND VGND VPWR VPWR _04865_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10965_ _05266_ net364 _05401_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12704_ clknet_leaf_120_clk _00162_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10896_ _04723_ _04724_ _04722_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__or3b_1
XFILLER_0_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12635_ clknet_leaf_142_clk _00093_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12566_ clknet_leaf_25_clk _01050_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11517_ _05304_ net631 _05706_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12497_ clknet_leaf_48_clk _00981_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 rvsingle.dp.rf.rf\[7\]\[17\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_888 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11448_ _05673_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11379_ _05635_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__clkbuf_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ clknet_leaf_133_clk _00576_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ clknet_leaf_10_clk _00507_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07610_ _01076_ _01071_ _01062_ _01145_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__a31o_1
X_08590_ _01694_ _03504_ _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07541_ _02452_ _02454_ _02461_ _01187_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07472_ _01675_ rvsingle.dp.rf.rf\[18\]\[6\] _01611_ _02392_ VGND VGND VPWR VPWR
+ _02393_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_159_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09211_ _04118_ _04119_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__a21oi_4
X_06423_ _01231_ _01339_ _01344_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09142_ _01250_ _04061_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__and2_1
X_06354_ _01099_ rvsingle.dp.rf.rf\[22\]\[29\] VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09073_ rvsingle.dp.rf.rf\[11\]\[26\] _01943_ _01451_ VGND VGND VPWR VPWR _03993_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06285_ _01207_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_170_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08024_ rvsingle.dp.rf.rf\[15\]\[0\] _01294_ _01243_ VGND VGND VPWR VPWR _02945_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold710 rvsingle.dp.rf.rf\[27\]\[29\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold721 rvsingle.dp.rf.rf\[23\]\[2\] VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold732 rvsingle.dp.rf.rf\[28\]\[19\] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold743 rvsingle.dp.rf.rf\[10\]\[25\] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold754 rvsingle.dp.rf.rf\[22\]\[22\] VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold765 rvsingle.dp.rf.rf\[24\]\[5\] VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 rvsingle.dp.rf.rf\[14\]\[12\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 rvsingle.dp.rf.rf\[25\]\[9\] VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 rvsingle.dp.rf.rf\[2\]\[1\] VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _04740_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__clkbuf_8
X_08926_ rvsingle.dp.rf.rf\[23\]\[25\] _03839_ _03840_ VGND VGND VPWR VPWR _03847_
+ sky130_fd_sc_hd__o21ai_1
X_08857_ _01842_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07808_ rvsingle.dp.rf.rf\[27\]\[3\] _01606_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__or2b_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _01426_ rvsingle.dp.rf.rf\[18\]\[15\] _01427_ VGND VGND VPWR VPWR _03709_
+ sky130_fd_sc_hd__o21a_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _02609_ _02658_ _01591_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__a21oi_2
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10750_ _05281_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09409_ _04260_ _04318_ _04321_ VGND VGND VPWR VPWR DataAdr[12] sky130_fd_sc_hd__o21ai_4
XFILLER_0_164_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10681_ _05243_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12420_ clknet_leaf_107_clk _00904_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12351_ _06127_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11302_ _05352_ rvsingle.dp.rf.rf\[15\]\[23\] _05591_ VGND VGND VPWR VPWR _05594_
+ sky130_fd_sc_hd__mux2_1
X_12282_ _05084_ _05835_ net215 VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11233_ _05354_ rvsingle.dp.rf.rf\[29\]\[24\] _05552_ VGND VGND VPWR VPWR _05556_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11164_ _05517_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10115_ _04713_ _04715_ _04138_ _04132_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__a22oi_1
X_11095_ _05460_ net191 _05181_ _05464_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__a22o_1
X_10046_ _01080_ _04612_ _04613_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__or3_2
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold70 rvsingle.dp.rf.rf\[15\]\[31\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 rvsingle.dp.rf.rf\[31\]\[31\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 rvsingle.dp.rf.rf\[7\]\[7\] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
X_11997_ _05965_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10948_ _05400_ net634 _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10879_ _05358_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12618_ clknet_leaf_83_clk _00076_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12549_ clknet_leaf_114_clk _01033_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ PC[20] _04582_ PC[21] VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__a21oi_1
X_06972_ rvsingle.dp.rf.rf\[21\]\[22\] _01865_ _01668_ _01892_ VGND VGND VPWR VPWR
+ _01893_ sky130_fd_sc_hd__o211ai_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _01567_ rvsingle.dp.rf.rf\[0\]\[14\] VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__nor2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _04533_ _04453_ _04535_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[14\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08642_ _02505_ _03537_ _03560_ _02375_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__a31oi_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08573_ rvsingle.dp.rf.rf\[11\]\[12\] _01901_ _03493_ VGND VGND VPWR VPWR _03494_
+ sky130_fd_sc_hd__o21ai_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07524_ rvsingle.dp.rf.rf\[7\]\[6\] _01687_ _01708_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07455_ _02375_ Instr[27] VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06406_ _01327_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__buf_8
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07386_ rvsingle.dp.rf.rf\[17\]\[7\] _02303_ _02285_ _02306_ VGND VGND VPWR VPWR
+ _02307_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09125_ _01614_ rvsingle.dp.rf.rf\[26\]\[26\] VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06337_ _01259_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__buf_4
XFILLER_0_161_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09056_ _03782_ _03968_ _03970_ _01117_ _03975_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__o311ai_4
X_06268_ _01190_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08007_ rvsingle.dp.rf.rf\[17\]\[0\] _01423_ _01454_ VGND VGND VPWR VPWR _02928_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_102_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold540 rvsingle.dp.rf.rf\[0\]\[1\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
X_06199_ rvsingle.dp.rf.rf\[8\]\[30\] rvsingle.dp.rf.rf\[9\]\[30\] rvsingle.dp.rf.rf\[10\]\[30\]
+ rvsingle.dp.rf.rf\[11\]\[30\] _01100_ _01120_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__mux4_1
Xhold551 rvsingle.dp.rf.rf\[0\]\[9\] VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 rvsingle.dp.rf.rf\[23\]\[17\] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 rvsingle.dp.rf.rf\[26\]\[17\] VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 rvsingle.dp.rf.rf\[10\]\[23\] VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 rvsingle.dp.rf.rf\[17\]\[11\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09958_ _04776_ _04468_ _04743_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__mux2_4
X_08909_ _03827_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__nand2_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _04713_ _04715_ _04118_ _04119_ _04129_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__a221oi_4
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _05901_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__clkbuf_8
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _05887_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__clkbuf_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _05187_ net447 _05298_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__mux2_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _05837_ net119 _05756_ _05841_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10733_ net9 _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10664_ _04917_ _04928_ _05057_ _04915_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_138_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12403_ clknet_leaf_35_clk _00887_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_100_clk _00811_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10595_ _04747_ rvsingle.dp.rf.rf\[22\]\[2\] _05194_ VGND VGND VPWR VPWR _05196_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ _06118_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12265_ _04823_ net435 _06073_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11216_ _05291_ rvsingle.dp.rf.rf\[29\]\[16\] _05541_ VGND VGND VPWR VPWR _05547_
+ sky130_fd_sc_hd__mux2_1
X_12196_ _04897_ net667 _06048_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11147_ _05476_ net658 _05499_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11078_ _04814_ _05145_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__nand2_1
X_10029_ _02909_ _02799_ _02910_ ReadData[20] _04715_ VGND VGND VPWR VPWR _04836_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07240_ rvsingle.dp.rf.rf\[8\]\[17\] rvsingle.dp.rf.rf\[9\]\[17\] _01241_ VGND VGND
+ VPWR VPWR _02161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07171_ rvsingle.dp.rf.rf\[27\]\[18\] _01943_ _02091_ VGND VGND VPWR VPWR _02092_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09812_ _04632_ _04635_ _04644_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__a21o_1
X_06955_ _01744_ rvsingle.dp.rf.rf\[24\]\[22\] VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__nor2_1
X_09743_ _04581_ _04582_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__or2_1
X_09674_ _04518_ _04519_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__xnor2_1
X_06886_ rvsingle.dp.rf.rf\[9\]\[23\] _01688_ _01689_ _01806_ VGND VGND VPWR VPWR
+ _01807_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_90_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _01545_ rvsingle.dp.rf.rf\[18\]\[12\] _02337_ _03545_ VGND VGND VPWR VPWR
+ _03546_ sky130_fd_sc_hd__o211ai_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08556_ _01463_ rvsingle.dp.rf.rf\[4\]\[13\] VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__nor2_1
X_07507_ _02427_ _01870_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08487_ _01658_ rvsingle.dp.rf.rf\[26\]\[13\] _01880_ _03407_ VGND VGND VPWR VPWR
+ _03408_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07438_ _01630_ rvsingle.dp.rf.rf\[20\]\[7\] VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07369_ _02288_ rvsingle.dp.rf.rf\[7\]\[7\] _01808_ _02289_ VGND VGND VPWR VPWR _02290_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09108_ rvsingle.dp.rf.rf\[11\]\[26\] _03778_ _04027_ VGND VGND VPWR VPWR _04028_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10380_ _04774_ net389 _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09039_ _01848_ rvsingle.dp.rf.rf\[2\]\[27\] _01612_ VGND VGND VPWR VPWR _03959_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12050_ _05173_ net476 _05983_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__mux2_1
Xhold370 rvsingle.dp.rf.rf\[25\]\[1\] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 rvsingle.dp.rf.rf\[8\]\[15\] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 rvsingle.dp.rf.rf\[23\]\[5\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _05432_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__clkbuf_1
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ clknet_leaf_23_clk _00410_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _05915_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__clkbuf_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _04978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12883_ clknet_leaf_34_clk _00341_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _05085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_232 _05499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 _01255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11834_ _05878_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__clkbuf_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _01695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_276 _01862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_287 _05004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11765_ _05837_ net101 _05745_ _05841_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__a22o_1
XANTENNA_298 _01513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10716_ _04870_ net365 _05257_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11696_ _05807_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10647_ _05224_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13366_ clknet_leaf_25_clk _00794_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10578_ _04892_ net294 _05151_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12317_ _06109_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13297_ clknet_leaf_59_clk _00755_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12248_ _04764_ rvsingle.dp.rf.rf\[5\]\[5\] _06074_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12179_ _05004_ _05348_ _06052_ net174 VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__a2bb2o_1
X_06740_ rvsingle.dp.rf.rf\[27\]\[20\] _01602_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__or2b_1
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06671_ _01152_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08410_ rvsingle.dp.rf.rf\[1\]\[9\] _01743_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09390_ _04303_ _04304_ _04136_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__nand3_4
XFILLER_0_58_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08341_ rvsingle.dp.rf.rf\[25\]\[8\] VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08272_ _03185_ _03187_ _01156_ _03192_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07223_ rvsingle.dp.rf.rf\[3\]\[17\] _01088_ _01626_ VGND VGND VPWR VPWR _02144_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07154_ rvsingle.dp.rf.rf\[8\]\[18\] rvsingle.dp.rf.rf\[9\]\[18\] rvsingle.dp.rf.rf\[10\]\[18\]
+ rvsingle.dp.rf.rf\[11\]\[18\] _01336_ _01200_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__mux4_2
XFILLER_0_15_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07085_ _02005_ rvsingle.dp.rf.rf\[4\]\[19\] _01530_ VGND VGND VPWR VPWR _02006_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07987_ _01081_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__clkbuf_4
X_06938_ _01855_ _01856_ _01512_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__a211oi_2
X_09726_ _04398_ _04563_ _04567_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[17\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06869_ rvsingle.dp.rf.rf\[17\]\[23\] _01558_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__and2b_1
X_09657_ PC[11] _04493_ _04497_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ rvsingle.dp.rf.rf\[7\]\[12\] _01650_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__and2b_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _04438_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ rvsingle.dp.rf.rf\[24\]\[13\] rvsingle.dp.rf.rf\[25\]\[13\] rvsingle.dp.rf.rf\[26\]\[13\]
+ rvsingle.dp.rf.rf\[27\]\[13\] _01468_ _01727_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__mux4_2
XFILLER_0_93_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11550_ _04754_ _05732_ _05733_ _05060_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__and4_1
XFILLER_0_147_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_987 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10501_ _05138_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11481_ _05330_ net686 _05684_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13220_ clknet_leaf_131_clk _00678_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10432_ _04879_ _04881_ _04880_ _04920_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__o31a_2
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13151_ clknet_leaf_0_clk _00609_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10363_ _05060_ _04970_ _05061_ net581 VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__a31o_1
X_12102_ _04785_ _04726_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__and2_1
X_13082_ clknet_leaf_6_clk _00540_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10294_ _05023_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__clkbuf_1
X_12033_ _05985_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ clknet_leaf_98_clk _00393_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12866_ clknet_leaf_140_clk _00324_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[23\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_75_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _05869_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ clknet_leaf_133_clk _00255_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11748_ _05724_ net808 _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11679_ _05798_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13418_ clknet_leaf_81_clk _00846_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13349_ clknet_leaf_79_clk rvsingle.dp.PCNext\[26\] _00026_ VGND VGND VPWR VPWR PC[26]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07910_ _02827_ _01716_ _02828_ _02830_ _02291_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__o311a_1
XFILLER_0_20_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08890_ rvsingle.dp.rf.rf\[24\]\[24\] rvsingle.dp.rf.rf\[25\]\[24\] rvsingle.dp.rf.rf\[26\]\[24\]
+ rvsingle.dp.rf.rf\[27\]\[24\] _01328_ _01455_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__mux4_1
X_07841_ _02756_ _01505_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__nand3_2
XFILLER_0_75_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07772_ _02690_ _02285_ _01206_ _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__a211o_1
X_09511_ _04391_ VGND VGND VPWR VPWR WriteData[4] sky130_fd_sc_hd__clkbuf_4
X_06723_ _01643_ rvsingle.dp.rf.rf\[30\]\[20\] VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09442_ DataAdr[3] _04345_ DataAdr[4] VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nor3_1
XFILLER_0_149_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06654_ _01497_ _01571_ _01572_ _01112_ _01574_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__o311ai_2
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09373_ _04284_ _04286_ _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06585_ _01505_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08324_ rvsingle.dp.rf.rf\[3\]\[8\] _02478_ _01523_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08255_ _03172_ _03173_ _03175_ _01600_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_15_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07206_ _01148_ rvsingle.dp.rf.rf\[8\]\[17\] VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__or2_1
X_08186_ rvsingle.dp.rf.rf\[9\]\[11\] _02379_ _01542_ _03106_ VGND VGND VPWR VPWR
+ _03107_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_144_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07137_ rvsingle.dp.rf.rf\[9\]\[18\] _01861_ _01759_ VGND VGND VPWR VPWR _02058_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07068_ _01744_ rvsingle.dp.rf.rf\[10\]\[19\] _01648_ _01988_ VGND VGND VPWR VPWR
+ _01989_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_100_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09709_ _04549_ _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__nor2_2
X_10981_ _05421_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12720_ clknet_leaf_52_clk _00178_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[18\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12651_ clknet_leaf_64_clk _00109_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[20\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11602_ _05713_ net299 _05729_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12582_ clknet_leaf_122_clk _00040_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11533_ _05719_ _05681_ _05720_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11464_ _05314_ _05681_ _05682_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13203_ clknet_leaf_48_clk _00661_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10415_ _04870_ net496 _05082_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11395_ _04739_ _05565_ _04738_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__or3b_2
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13134_ clknet_leaf_71_clk _00592_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10346_ _05050_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__clkbuf_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ clknet_leaf_89_clk _00523_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10277_ _04886_ rvsingle.dp.rf.rf\[27\]\[27\] _05001_ VGND VGND VPWR VPWR _05013_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12016_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__buf_6
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap2 _03454_ VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__buf_2
X_12918_ clknet_leaf_32_clk _00376_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12849_ clknet_leaf_48_clk _00307_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06370_ _01210_ _01291_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08040_ _01315_ _02949_ _02960_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09991_ _02909_ _02799_ _02910_ ReadData[14] _04715_ VGND VGND VPWR VPWR _04804_
+ sky130_fd_sc_hd__o311a_1
X_08942_ _03778_ rvsingle.dp.rf.rf\[7\]\[25\] _01106_ _03862_ VGND VGND VPWR VPWR
+ _03863_ sky130_fd_sc_hd__o211ai_1
X_08873_ _03782_ _03793_ _01506_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07824_ _02732_ _02744_ _01145_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__nand3_2
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07755_ _02163_ rvsingle.dp.rf.rf\[12\]\[3\] VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06706_ _01256_ rvsingle.dp.rf.rf\[4\]\[20\] VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07686_ _02599_ _02606_ _01187_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__nand3_1
XFILLER_0_149_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09425_ _02803_ _02851_ _02861_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__o21ai_1
X_06637_ _01557_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__buf_6
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09356_ _04220_ _04223_ _04271_ _04136_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__o211ai_1
X_06568_ _01103_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08307_ _03124_ _03139_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nand2_1
X_09287_ _01583_ _01589_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__nand3_1
X_06499_ _01419_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__buf_8
X_08238_ rvsingle.dp.rf.rf\[15\]\[10\] _01901_ _03158_ VGND VGND VPWR VPWR _03159_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08169_ _01381_ rvsingle.dp.rf.rf\[6\]\[11\] VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10200_ _04909_ _04913_ _04923_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11180_ _05314_ _05525_ _05526_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__a21oi_1
X_10131_ _04924_ _04925_ net24 VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10062_ _04864_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10964_ _05410_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12703_ clknet_leaf_131_clk _00161_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10895_ _05314_ _05368_ _05369_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12634_ clknet_leaf_3_clk _00092_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12565_ clknet_leaf_64_clk _01049_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11516_ _05710_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12496_ clknet_leaf_70_clk _00980_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11447_ _05304_ rvsingle.dp.rf.rf\[13\]\[25\] _05668_ VGND VGND VPWR VPWR _05673_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11378_ _05407_ net512 _05629_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10329_ _05041_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__clkbuf_1
X_13117_ clknet_leaf_145_clk _00575_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ clknet_leaf_10_clk _00506_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07540_ _01229_ _02455_ _02460_ _02447_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07471_ rvsingle.dp.rf.rf\[19\]\[6\] _01096_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06422_ _01341_ _01231_ _01343_ _01222_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__a31o_1
X_09210_ _04128_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09141_ _01182_ _01186_ _01249_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__a21o_1
X_06353_ rvsingle.dp.rf.rf\[20\]\[29\] rvsingle.dp.rf.rf\[21\]\[29\] _01139_ VGND
+ VGND VPWR VPWR _01276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09072_ _03989_ _01310_ _01209_ _03991_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_142_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06284_ _01206_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__buf_6
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08023_ _01328_ rvsingle.dp.rf.rf\[14\]\[0\] VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold700 rvsingle.dp.rf.rf\[30\]\[20\] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold711 rvsingle.dp.rf.rf\[22\]\[16\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold722 rvsingle.dp.rf.rf\[27\]\[26\] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold733 rvsingle.dp.rf.rf\[26\]\[13\] VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold744 rvsingle.dp.rf.rf\[15\]\[15\] VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 rvsingle.dp.rf.rf\[28\]\[17\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 rvsingle.dp.rf.rf\[29\]\[1\] VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 rvsingle.dp.rf.rf\[8\]\[8\] VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold788 rvsingle.dp.rf.rf\[15\]\[20\] VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 rvsingle.dp.rf.rf\[7\]\[2\] VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08925_ _01257_ rvsingle.dp.rf.rf\[22\]\[25\] VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__nor2_1
X_08856_ _03776_ _01497_ _01565_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07807_ rvsingle.dp.rf.rf\[25\]\[3\] _01779_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__and2b_1
XFILLER_0_169_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08787_ rvsingle.dp.rf.rf\[17\]\[15\] _01424_ _02285_ _03707_ VGND VGND VPWR VPWR
+ _03708_ sky130_fd_sc_hd__o211ai_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _01065_ _01074_ _02609_ _02658_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__o211a_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07669_ _02587_ _01689_ _01702_ _02589_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09408_ _03513_ _04319_ _03564_ _04320_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__o211ai_2
X_10680_ _04778_ net683 _05235_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09339_ _02151_ _04254_ _04143_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12350_ _04876_ net268 _06121_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11301_ _05593_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__clkbuf_1
X_12281_ _06074_ net134 _05182_ _05832_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11232_ _05555_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11163_ _05304_ net335 _05511_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10114_ _04879_ _04880_ _04881_ ReadData[31] _04715_ VGND VGND VPWR VPWR _04910_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11094_ _05480_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__clkbuf_1
X_10045_ _04751_ _04210_ _04849_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold60 rvsingle.dp.rf.rf\[11\]\[6\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 rvsingle.dp.rf.rf\[14\]\[31\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold82 rvsingle.dp.rf.rf\[5\]\[15\] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 rvsingle.dp.rf.rf\[11\]\[10\] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
X_11996_ _05132_ net375 _05960_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10947_ _05372_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__buf_8
XFILLER_0_58_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10878_ _05307_ rvsingle.dp.rf.rf\[1\]\[27\] _05319_ VGND VGND VPWR VPWR _05358_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12617_ clknet_leaf_95_clk _00075_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_979 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12548_ clknet_leaf_107_clk _01032_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12479_ clknet_leaf_1_clk _00963_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_2 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _01675_ rvsingle.dp.rf.rf\[20\]\[22\] VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__or2_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _03625_ _02527_ _03630_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__nand3_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _04454_ _04455_ _04534_ _04459_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__o211ai_1
X_08641_ _01537_ _01171_ _01183_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__o211ai_4
X_08572_ _02450_ rvsingle.dp.rf.rf\[10\]\[12\] _01427_ VGND VGND VPWR VPWR _03493_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07523_ _01707_ rvsingle.dp.rf.rf\[6\]\[6\] VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07454_ net822 VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06405_ Instr[15] VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07385_ _01462_ rvsingle.dp.rf.rf\[16\]\[7\] VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06336_ _01258_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__buf_6
X_09124_ _01488_ rvsingle.dp.rf.rf\[25\]\[26\] _04043_ VGND VGND VPWR VPWR _04044_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09055_ _03972_ _01512_ _03974_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__nand3_1
XFILLER_0_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06267_ Instr[15] VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08006_ _02450_ rvsingle.dp.rf.rf\[16\]\[0\] VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__nor2_1
Xhold530 rvsingle.dp.rf.rf\[8\]\[14\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06198_ _01114_ _01121_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__nor2_1
Xhold541 rvsingle.dp.rf.rf\[11\]\[18\] VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold552 rvsingle.dp.rf.rf\[10\]\[15\] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 rvsingle.dp.rf.rf\[19\]\[1\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 rvsingle.dp.rf.rf\[30\]\[22\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 rvsingle.dp.rf.rf\[8\]\[5\] VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 rvsingle.dp.rf.rf\[5\]\[23\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ DataAdr[8] ReadData[8] _04751_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__mux2_1
X_08908_ _03828_ _03803_ _03825_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__o21bai_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _04245_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__clkbuf_4
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _02015_ _02016_ _02098_ _02100_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__nand4_1
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _04852_ net635 _05885_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__mux2_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _05310_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11781_ _05850_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__clkbuf_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10732_ _04917_ _04920_ _04922_ _04916_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__and4b_2
XFILLER_0_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10663_ _04719_ _05232_ _05233_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12402_ clknet_leaf_41_clk _00886_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10594_ _05195_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__clkbuf_1
X_13382_ clknet_leaf_122_clk _00810_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12333_ _05173_ net760 _06110_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12264_ _06082_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11215_ _05546_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__clkbuf_1
X_12195_ _06063_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11146_ _05508_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11077_ _05169_ _05471_ _05463_ net158 VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10028_ _04835_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11979_ _05956_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07170_ _01242_ rvsingle.dp.rf.rf\[26\]\[18\] _01471_ VGND VGND VPWR VPWR _02091_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_120_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09811_ _04632_ _04635_ _04644_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nand3_1
X_09742_ PC[17] PC[18] PC[19] _04554_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__and4_1
X_06954_ _01871_ _01872_ _01112_ _01874_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09673_ _04511_ _04504_ _04509_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__o21ba_1
X_06885_ _01707_ rvsingle.dp.rf.rf\[8\]\[23\] VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ rvsingle.dp.rf.rf\[19\]\[12\] _02627_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08555_ rvsingle.dp.rf.rf\[7\]\[13\] _02303_ _01199_ VGND VGND VPWR VPWR _03476_
+ sky130_fd_sc_hd__o21ai_2
X_07506_ _01139_ _01962_ _02402_ _02426_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__o211ai_4
X_08486_ rvsingle.dp.rf.rf\[27\]\[13\] _01381_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__or2b_1
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07437_ _02348_ _02352_ _01505_ _02357_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_9_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07368_ _01828_ rvsingle.dp.rf.rf\[6\]\[7\] VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09107_ _01848_ rvsingle.dp.rf.rf\[10\]\[26\] _01612_ VGND VGND VPWR VPWR _04027_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06319_ _01241_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_111_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_111_clk sky130_fd_sc_hd__clkbuf_16
X_07299_ rvsingle.dp.rf.rf\[23\]\[16\] _01513_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__or2b_1
XFILLER_0_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09038_ _03857_ rvsingle.dp.rf.rf\[1\]\[27\] _03957_ VGND VGND VPWR VPWR _03958_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold360 rvsingle.dp.rf.rf\[6\]\[16\] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 rvsingle.dp.rf.rf\[25\]\[30\] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 rvsingle.dp.rf.rf\[26\]\[27\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 rvsingle.dp.rf.rf\[28\]\[2\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _05334_ net815 _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__mux2_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ clknet_leaf_9_clk _00409_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _04795_ net526 _05913_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _04384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12882_ clknet_leaf_41_clk _00340_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _04978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _05085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11833_ _05391_ net246 _05874_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__mux2_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 rvsingle.dp.rf.rf\[24\]\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _01426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_266 _01726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _05844_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_288 _05004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_299 _01603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _05261_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _05744_ rvsingle.dp.rf.rf\[10\]\[11\] _05806_ VGND VGND VPWR VPWR _05807_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10646_ _04870_ net747 _05219_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_102_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13365_ clknet_leaf_64_clk _00793_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10577_ _04886_ _05183_ _05146_ _05184_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12316_ _04785_ net525 _06099_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13296_ clknet_leaf_67_clk _00754_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12247_ _06077_ net181 _05465_ _05832_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12178_ net20 _06049_ _05347_ _05766_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__a22o_1
X_11129_ _05330_ rvsingle.dp.rf.rf\[16\]\[8\] _05499_ VGND VGND VPWR VPWR _05500_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06670_ _01485_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__buf_4
XFILLER_0_114_1002 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_974 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08340_ _01605_ _03256_ _03257_ _01511_ _03260_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__o311a_1
XFILLER_0_171_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08271_ _01605_ _03188_ _03189_ _01511_ _03191_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07222_ _01666_ rvsingle.dp.rf.rf\[2\]\[17\] VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07153_ _01915_ _02069_ _02073_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_144_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07084_ _01124_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__buf_6
XFILLER_0_113_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07986_ _01592_ _02885_ _02906_ _01178_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__a31oi_4
X_09725_ _04422_ _04423_ _04566_ _04427_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__o211a_1
X_06937_ _01848_ rvsingle.dp.rf.rf\[2\]\[22\] _01612_ _01857_ VGND VGND VPWR VPWR
+ _01858_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09656_ _04499_ _04453_ _04503_ VGND VGND VPWR VPWR rvsingle.dp.PCNext\[11\] sky130_fd_sc_hd__o21ai_1
X_06868_ _01137_ rvsingle.dp.rf.rf\[16\]\[23\] _01611_ VGND VGND VPWR VPWR _01789_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _01558_ rvsingle.dp.rf.rf\[6\]\[12\] _01777_ VGND VGND VPWR VPWR _03528_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ Instr[25] _04429_ _04439_ _04419_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__o22a_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ _01715_ _01717_ _01703_ _01719_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__a211oi_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _01207_ _03458_ _02447_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08469_ rvsingle.dp.rf.rf\[20\]\[9\] rvsingle.dp.rf.rf\[21\]\[9\] rvsingle.dp.rf.rf\[22\]\[9\]
+ rvsingle.dp.rf.rf\[23\]\[9\] _01328_ _01455_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10500_ _04898_ net341 _05126_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11480_ _05691_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10431_ _05097_ _04924_ _04970_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13150_ clknet_leaf_0_clk _00608_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10362_ _05057_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__buf_4
X_12101_ _06020_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__clkbuf_1
X_10293_ _04736_ net762 _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__mux2_1
X_13081_ clknet_leaf_9_clk _00539_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12032_ _05740_ net777 _05983_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__mux2_1
Xhold190 rvsingle.dp.rf.rf\[7\]\[25\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ clknet_leaf_114_clk _00392_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ clknet_leaf_140_clk _00323_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _05496_ net779 _05863_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__mux2_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ clknet_leaf_149_clk _00254_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11747_ _05836_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__buf_8
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11678_ _05531_ rvsingle.dp.rf.rf\[10\]\[3\] _05795_ VGND VGND VPWR VPWR _05798_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13417_ clknet_leaf_94_clk _00845_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10629_ _04824_ net369 _05205_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13348_ clknet_leaf_78_clk rvsingle.dp.PCNext\[25\] _00025_ VGND VGND VPWR VPWR PC[25]
+ sky130_fd_sc_hd__dfrtp_4
X_13279_ clknet_leaf_135_clk _00737_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07840_ _02758_ _02410_ _02760_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07771_ _01423_ rvsingle.dp.rf.rf\[31\]\[3\] _02691_ VGND VGND VPWR VPWR _02692_
+ sky130_fd_sc_hd__o21a_1
X_09510_ _04377_ _02504_ _02529_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__and3_4
X_06722_ _01642_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09441_ _04346_ _04135_ _04347_ _04348_ VGND VGND VPWR VPWR DataAdr[4] sky130_fd_sc_hd__a31o_4
X_06653_ _01540_ rvsingle.dp.rf.rf\[5\]\[21\] _01573_ VGND VGND VPWR VPWR _01574_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09372_ _04059_ _04180_ _04137_ _04287_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__o211ai_4
X_06584_ _01115_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__buf_8
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08323_ _01137_ rvsingle.dp.rf.rf\[2\]\[8\] VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08254_ _01595_ rvsingle.dp.rf.rf\[8\]\[10\] _03174_ _02485_ VGND VGND VPWR VPWR
+ _03175_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07205_ _02113_ _02125_ _01682_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__nand3_4
X_08185_ _01096_ rvsingle.dp.rf.rf\[8\]\[11\] VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07136_ _01559_ rvsingle.dp.rf.rf\[8\]\[18\] VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07067_ rvsingle.dp.rf.rf\[11\]\[19\] _01753_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__or2b_1
XFILLER_0_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07969_ _02886_ _02887_ _01617_ _02889_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09708_ _04527_ _04528_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__a21oi_2
X_10980_ _05322_ net689 _05419_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09639_ _04481_ _04482_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__nand2_1
X_12650_ clknet_leaf_82_clk _00108_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11601_ _05761_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12581_ clknet_leaf_123_clk _00039_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11532_ _05364_ _05365_ _05681_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11463_ net136 _05681_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__nor2_1
X_13202_ clknet_leaf_53_clk _00660_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10414_ _05088_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11394_ _05314_ _05643_ _05644_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13133_ clknet_leaf_45_clk _00591_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10345_ _04877_ net405 _05044_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ clknet_leaf_103_clk _00522_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _05012_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_1
X_12015_ _04737_ _04919_ _04733_ _05149_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__or4_4
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12917_ clknet_leaf_37_clk _00375_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12848_ clknet_leaf_53_clk _00306_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ clknet_leaf_86_clk _00237_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09990_ _04803_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
X_08941_ _01643_ rvsingle.dp.rf.rf\[6\]\[25\] VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08872_ rvsingle.dp.rf.rf\[8\]\[24\] rvsingle.dp.rf.rf\[9\]\[24\] rvsingle.dp.rf.rf\[10\]\[24\]
+ rvsingle.dp.rf.rf\[11\]\[24\] _01518_ _01626_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07823_ _02735_ _02738_ _02364_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07754_ rvsingle.dp.rf.rf\[8\]\[3\] rvsingle.dp.rf.rf\[9\]\[3\] rvsingle.dp.rf.rf\[10\]\[3\]
+ rvsingle.dp.rf.rf\[11\]\[3\] _02176_ _01696_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__mux4_1
XFILLER_0_168_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06705_ _01611_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07685_ _01422_ _02600_ _02605_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_91_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
X_09424_ _02751_ _02856_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__and2_1
X_06636_ _01095_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09355_ _03738_ _03739_ _03573_ _04259_ _04162_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__o221ai_1
X_06567_ _01487_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08306_ _03222_ _03223_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__nand3_4
XFILLER_0_145_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09286_ _04146_ _04167_ _01739_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06498_ _01190_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08237_ _01903_ rvsingle.dp.rf.rf\[14\]\[10\] _01243_ VGND VGND VPWR VPWR _03158_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08168_ rvsingle.dp.rf.rf\[5\]\[11\] _01613_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__and2b_1
X_07119_ _01634_ _02034_ _02039_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__nand3_1
X_08099_ _01602_ rvsingle.dp.rf.rf\[20\]\[1\] VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10130_ _04722_ _04723_ _04921_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__and3_2
XFILLER_0_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10061_ _04863_ net420 _04847_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10963_ _05359_ net340 _05401_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_16
X_12702_ clknet_leaf_133_clk _00160_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10894_ net115 _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12633_ clknet_leaf_8_clk _00091_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12564_ clknet_leaf_21_clk _01048_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11515_ _05354_ rvsingle.dp.rf.rf\[12\]\[24\] _05706_ VGND VGND VPWR VPWR _05710_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12495_ clknet_leaf_39_clk _00979_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11446_ _05672_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11377_ _05634_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13116_ clknet_leaf_13_clk _00574_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10328_ _04828_ net418 _05033_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__mux2_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ clknet_leaf_11_clk _00505_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10259_ _04505_ _01071_ _01062_ _04975_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__a31o_4
XFILLER_0_89_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_73_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07470_ rvsingle.dp.rf.rf\[17\]\[6\] _01594_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__and2b_1
X_06421_ rvsingle.dp.rf.rf\[23\]\[29\] _01297_ _01342_ VGND VGND VPWR VPWR _01343_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09140_ _01348_ _01410_ _01415_ _04059_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__o22ai_4
X_06352_ _01113_ _01274_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09071_ _01297_ rvsingle.dp.rf.rf\[7\]\[26\] _01201_ _03990_ VGND VGND VPWR VPWR
+ _03991_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06283_ Instr[17] VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08022_ _02873_ _01707_ _02942_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold701 rvsingle.dp.rf.rf\[14\]\[1\] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold712 rvsingle.dp.rf.rf\[18\]\[11\] VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 rvsingle.dp.rf.rf\[13\]\[16\] VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold734 rvsingle.dp.rf.rf\[6\]\[5\] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold745 rvsingle.dp.rf.rf\[22\]\[11\] VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 rvsingle.dp.rf.rf\[21\]\[26\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 rvsingle.dp.rf.rf\[9\]\[11\] VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 rvsingle.dp.rf.rf\[23\]\[7\] VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _04788_ _04502_ _04743_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__mux2_4
Xhold789 rvsingle.dp.rf.rf\[26\]\[6\] VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ rvsingle.dp.rf.rf\[21\]\[25\] _01643_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__and2b_1
X_08855_ rvsingle.dp.rf.rf\[20\]\[24\] rvsingle.dp.rf.rf\[21\]\[24\] _01780_ VGND
+ VGND VPWR VPWR _03776_ sky130_fd_sc_hd__mux2_1
X_07806_ _01125_ rvsingle.dp.rf.rf\[24\]\[3\] VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__nor2_1
X_08786_ _02440_ rvsingle.dp.rf.rf\[16\]\[15\] VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__or2_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _02633_ _01083_ _02505_ _02657_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__nand4_2
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_64_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07668_ _02271_ rvsingle.dp.rf.rf\[11\]\[5\] _01300_ _02588_ VGND VGND VPWR VPWR
+ _02589_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09407_ Instr[13] Instr[14] _04141_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__and3_2
X_06619_ _01539_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07599_ _01595_ rvsingle.dp.rf.rf\[28\]\[4\] _02519_ _02485_ VGND VGND VPWR VPWR
+ _02520_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_47_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09338_ _01185_ _02261_ _02152_ _02181_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09269_ _01348_ _01410_ _01415_ _04059_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11300_ _05300_ rvsingle.dp.rf.rf\[15\]\[22\] _05591_ VGND VGND VPWR VPWR _05593_
+ sky130_fd_sc_hd__mux2_1
X_12280_ _06089_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11231_ _05352_ rvsingle.dp.rf.rf\[29\]\[23\] _05552_ VGND VGND VPWR VPWR _05555_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11162_ _05490_ net197 _05133_ _05501_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10113_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11093_ _05354_ rvsingle.dp.rf.rf\[17\]\[24\] _05469_ VGND VGND VPWR VPWR _05480_
+ sky130_fd_sc_hd__mux2_1
X_10044_ _02909_ _02799_ _02910_ ReadData[22] _04245_ VGND VGND VPWR VPWR _04849_
+ sky130_fd_sc_hd__o311a_1
Xhold50 rvsingle.dp.rf.rf\[9\]\[10\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 rvsingle.dp.rf.rf\[0\]\[31\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 rvsingle.dp.rf.rf\[19\]\[7\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 rvsingle.dp.rf.rf\[5\]\[14\] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold94 rvsingle.dp.rf.rf\[9\]\[19\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
X_11995_ _05964_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_55_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10946_ _04845_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__buf_2
XFILLER_0_86_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10877_ _05357_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12616_ clknet_leaf_106_clk _00074_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12547_ clknet_leaf_127_clk _01031_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12478_ clknet_leaf_150_clk _00962_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_3 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11429_ _05663_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06970_ rvsingle.dp.rf.rf\[23\]\[22\] _01865_ _01626_ VGND VGND VPWR VPWR _01891_
+ sky130_fd_sc_hd__o21ai_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08640_ _02505_ _03537_ _03560_ _01177_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08571_ rvsingle.dp.rf.rf\[9\]\[12\] _01295_ _02285_ VGND VGND VPWR VPWR _03492_
+ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_46_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07522_ rvsingle.dp.rf.rf\[5\]\[6\] _01687_ _02268_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07453_ _02317_ _02373_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06404_ rvsingle.dp.rf.rf\[28\]\[29\] rvsingle.dp.rf.rf\[29\]\[29\] _01194_ VGND
+ VGND VPWR VPWR _01326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07384_ _02303_ rvsingle.dp.rf.rf\[19\]\[7\] _01953_ _02304_ VGND VGND VPWR VPWR
+ _02305_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09123_ _01614_ rvsingle.dp.rf.rf\[24\]\[26\] VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06335_ Instr[21] VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__buf_8
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09054_ rvsingle.dp.rf.rf\[15\]\[27\] _03857_ _03973_ VGND VGND VPWR VPWR _03974_
+ sky130_fd_sc_hd__o21ai_1
X_06266_ _01188_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08005_ _02273_ _02920_ _02925_ _01446_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_170_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold520 rvsingle.dp.rf.rf\[6\]\[19\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06197_ rvsingle.dp.rf.rf\[0\]\[30\] rvsingle.dp.rf.rf\[1\]\[30\] rvsingle.dp.rf.rf\[2\]\[30\]
+ rvsingle.dp.rf.rf\[3\]\[30\] _01100_ _01120_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__mux4_1
Xhold531 rvsingle.dp.rf.rf\[0\]\[14\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 rvsingle.dp.rf.rf\[6\]\[4\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold553 rvsingle.dp.rf.rf\[6\]\[30\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 rvsingle.dp.rf.rf\[11\]\[30\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold575 rvsingle.dp.rf.rf\[22\]\[7\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold586 rvsingle.dp.rf.rf\[25\]\[4\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 rvsingle.dp.rf.rf\[26\]\[16\] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09956_ _04775_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
X_08907_ _01961_ Instr[31] _01184_ _03802_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__a211oi_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ ReadData[0] _01080_ _04121_ _04713_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__and4b_1
XFILLER_0_99_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _03064_ _03736_ _03758_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a21oi_4
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08769_ _01545_ rvsingle.dp.rf.rf\[4\]\[15\] VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_37_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _05266_ net461 _05298_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__mux2_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _04845_ net310 _05845_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__mux2_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10731_ _05269_ _05232_ _05270_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10662_ net127 _05232_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_982 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12401_ clknet_leaf_49_clk _00885_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13381_ clknet_leaf_123_clk _00809_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10593_ _04736_ net735 _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12332_ _06117_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12263_ _05344_ net232 _06074_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__mux2_1
X_11214_ _05212_ rvsingle.dp.rf.rf\[29\]\[15\] _05541_ VGND VGND VPWR VPWR _05546_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12194_ _05763_ net324 _06048_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11145_ _05291_ net522 _05499_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11076_ _05473_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__clkbuf_1
X_10027_ _04834_ net615 _04791_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
X_11978_ _04813_ net655 _05949_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10929_ _05390_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09810_ _04617_ PC[25] VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__xnor2_2
X_09741_ PC[17] PC[18] _04554_ PC[19] VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__a31oi_1
X_06953_ rvsingle.dp.rf.rf\[29\]\[22\] _01861_ _01759_ _01873_ VGND VGND VPWR VPWR
+ _01874_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09672_ _04516_ _04517_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__or2b_1
X_06884_ rvsingle.dp.rf.rf\[12\]\[23\] rvsingle.dp.rf.rf\[13\]\[23\] rvsingle.dp.rf.rf\[14\]\[23\]
+ rvsingle.dp.rf.rf\[15\]\[23\] _01417_ _01301_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08623_ rvsingle.dp.rf.rf\[17\]\[12\] _03258_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_19_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _01463_ rvsingle.dp.rf.rf\[6\]\[13\] VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07505_ _01377_ _02414_ _02425_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__nand3_4
XFILLER_0_49_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08485_ _03313_ _03317_ _03399_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__nand4_2
X_07436_ _02320_ _02353_ _02354_ _02323_ _02356_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07367_ _01294_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__buf_6
XFILLER_0_73_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09106_ rvsingle.dp.rf.rf\[9\]\[26\] _03857_ _01856_ VGND VGND VPWR VPWR _04026_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06318_ _01240_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07298_ _01269_ rvsingle.dp.rf.rf\[20\]\[16\] _02218_ _01497_ VGND VGND VPWR VPWR
+ _02219_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_131_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09037_ _01848_ rvsingle.dp.rf.rf\[0\]\[27\] _01605_ VGND VGND VPWR VPWR _03957_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06249_ Instr[17] VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold350 rvsingle.dp.rf.rf\[27\]\[1\] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 rvsingle.dp.rf.rf\[16\]\[30\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 rvsingle.dp.rf.rf\[9\]\[15\] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 rvsingle.dp.rf.rf\[1\]\[7\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 rvsingle.dp.rf.rf\[28\]\[27\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09939_ _04761_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ clknet_leaf_31_clk _00408_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _05914_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__clkbuf_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ clknet_leaf_42_clk _00339_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[15\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _04388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _05000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ _05877_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__clkbuf_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 _05775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_245 rvsingle.dp.rf.rf\[24\]\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _01437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_267 _01777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 _02150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _05385_ net588 _05837_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 _05004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _04863_ net411 _05257_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__mux2_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11694_ _05794_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__buf_6
XFILLER_0_165_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10645_ _05223_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13364_ clknet_4_12_0_clk _00792_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10576_ _05145_ _05146_ _03924_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12315_ _06108_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__clkbuf_1
X_13295_ clknet_leaf_44_clk _00753_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12246_ _06077_ net45 _05156_ _05841_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12177_ net103 _06049_ _05346_ _05766_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__a22o_1
X_11128_ _05489_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__buf_8
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11059_ net198 _05460_ _05465_ _05464_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_986 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08270_ rvsingle.dp.rf.rf\[7\]\[10\] _02481_ _03190_ VGND VGND VPWR VPWR _03191_
+ sky130_fd_sc_hd__o21ai_1
X_07221_ _02138_ _02139_ _01503_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07152_ _02070_ _01717_ _01722_ _02072_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07083_ rvsingle.dp.rf.rf\[7\]\[19\] _01675_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07985_ _02890_ _02895_ _02900_ _02905_ _01682_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__o221ai_4
X_09724_ _04564_ _04565_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__nand2_1
X_06936_ rvsingle.dp.rf.rf\[3\]\[22\] _01658_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__or2b_1
XFILLER_0_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09655_ _04454_ _04455_ _04502_ _04459_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__o211ai_1
X_06867_ _01776_ _01782_ _01526_ _01787_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__o211ai_1
X_08606_ _03525_ _01256_ _01531_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09586_ Instr[25] _04429_ _02532_ PC[4] VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__a22o_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ _01688_ rvsingle.dp.rf.rf\[19\]\[20\] _01456_ _01718_ VGND VGND VPWR VPWR
+ _01719_ sky130_fd_sc_hd__o211a_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ rvsingle.dp.rf.rf\[20\]\[13\] rvsingle.dp.rf.rf\[21\]\[13\] rvsingle.dp.rf.rf\[22\]\[13\]
+ rvsingle.dp.rf.rf\[23\]\[13\] _01328_ _01470_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08468_ _02093_ _03383_ _03388_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07419_ _02117_ rvsingle.dp.rf.rf\[4\]\[7\] VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08399_ rvsingle.dp.rf.rf\[9\]\[9\] _01607_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10430_ _04720_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10361_ _04720_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__clkbuf_8
X_12100_ _04781_ net551 _06019_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13080_ clknet_leaf_22_clk _00538_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10292_ _05021_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__buf_8
XFILLER_0_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12031_ _05984_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__clkbuf_1
Xhold180 rvsingle.dp.rf.rf\[0\]\[26\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold191 rvsingle.dp.rf.rf\[17\]\[25\] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ clknet_leaf_108_clk _00391_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ clknet_leaf_116_clk _00322_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _05868_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12795_ clknet_leaf_142_clk _00253_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[17\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11746_ _04505_ _01071_ _01062_ _05417_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__a311o_4
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11677_ _05797_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13416_ clknet_leaf_106_clk _00844_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[30\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_10628_ _05214_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13347_ clknet_leaf_78_clk rvsingle.dp.PCNext\[24\] _00024_ VGND VGND VPWR VPWR PC[24]
+ sky130_fd_sc_hd__dfrtp_4
X_10559_ _04834_ _05145_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13278_ clknet_leaf_146_clk _00736_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12229_ _06069_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__inv_2
X_07770_ _01425_ rvsingle.dp.rf.rf\[30\]\[3\] _01197_ VGND VGND VPWR VPWR _02691_
+ sky130_fd_sc_hd__o21a_1
X_06721_ _01606_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09440_ _02570_ _02534_ _02572_ _04142_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__o211a_1
X_06652_ _01499_ rvsingle.dp.rf.rf\[4\]\[21\] _01259_ VGND VGND VPWR VPWR _01573_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09371_ _04059_ _04180_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06583_ _01497_ _01500_ _01501_ _01503_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08322_ _03237_ _03242_ _02527_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__nand3_2
XFILLER_0_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08253_ rvsingle.dp.rf.rf\[9\]\[10\] _01594_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__or2b_1
XFILLER_0_144_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_894 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07204_ _02116_ _02119_ _01634_ _02124_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_144_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08184_ rvsingle.dp.rf.rf\[11\]\[11\] _01860_ _01880_ VGND VGND VPWR VPWR _03105_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07135_ _02052_ _02053_ _01112_ _02055_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_132_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07066_ rvsingle.dp.rf.rf\[9\]\[19\] _01382_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07968_ rvsingle.dp.rf.rf\[31\]\[0\] _01646_ _02888_ VGND VGND VPWR VPWR _02889_
+ sky130_fd_sc_hd__o21ai_1
X_06919_ _01836_ _01839_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__nand2_2
X_09707_ _04530_ _04539_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__or2_1
X_07899_ _01691_ rvsingle.dp.rf.rf\[6\]\[2\] VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09638_ _04481_ _04482_ _04484_ _04486_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_167_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09569_ _04397_ PC[3] PC[4] VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11600_ _05407_ net617 _05729_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12580_ clknet_leaf_123_clk _00038_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11531_ net38 VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11462_ _04916_ _04918_ _04920_ _04922_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__and4b_2
XFILLER_0_163_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13201_ clknet_leaf_55_clk _00659_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10413_ _04863_ net308 _05082_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11393_ net178 _05643_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13132_ clknet_leaf_48_clk _00590_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[23\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10344_ _05049_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ clknet_leaf_97_clk _00521_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10275_ _04877_ net722 _05001_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__mux2_1
X_12014_ _05721_ _05973_ _05974_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap4 _01177_ VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__buf_4
X_12916_ clknet_leaf_61_clk _00374_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[14\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ clknet_leaf_37_clk _00305_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[29\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ clknet_leaf_81_clk _00236_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[31\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11729_ _05824_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08940_ _03856_ _03858_ _03859_ _03860_ _02236_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__o221a_1
X_08871_ _02236_ _03791_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__nor2_1
X_07822_ _01777_ _02739_ _02740_ _01599_ _02742_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07753_ _01207_ _02673_ _02447_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__o21ai_1
X_06704_ rvsingle.dp.rf.rf\[5\]\[20\] VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__inv_2
X_07684_ _01460_ _02602_ _02604_ _01215_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_149_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09423_ _02854_ _02750_ _02855_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__o21ai_1
X_06635_ _01548_ _01555_ _01506_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__nand3_1
XFILLER_0_149_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09354_ _04121_ _04122_ _03645_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06566_ _01086_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08305_ _03224_ _03225_ _01584_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09285_ _01180_ _03978_ _03981_ _04200_ _04143_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__o221ai_4
X_06497_ rvsingle.dp.rf.rf\[24\]\[21\] rvsingle.dp.rf.rf\[25\]\[21\] rvsingle.dp.rf.rf\[26\]\[21\]
+ rvsingle.dp.rf.rf\[27\]\[21\] _01417_ _01301_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08236_ rvsingle.dp.rf.rf\[13\]\[10\] _01901_ _02285_ _03156_ VGND VGND VPWR VPWR
+ _03157_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_145_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08167_ _01097_ rvsingle.dp.rf.rf\[4\]\[11\] VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07118_ _01260_ _02035_ _02036_ _01503_ _02038_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08098_ _03002_ _03007_ _01376_ _03018_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_100_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07049_ _01148_ rvsingle.dp.rf.rf\[22\]\[19\] _01611_ VGND VGND VPWR VPWR _01970_
+ sky130_fd_sc_hd__o21a_1
X_10060_ _04862_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10962_ _05409_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12701_ clknet_leaf_136_clk _00159_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10893_ _04721_ _04728_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__and3_2
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12632_ clknet_leaf_33_clk _00090_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[21\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12563_ clknet_4_8_0_clk _01047_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11514_ _05709_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12494_ clknet_leaf_67_clk _00978_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[25\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11445_ _05354_ rvsingle.dp.rf.rf\[13\]\[24\] _05668_ VGND VGND VPWR VPWR _05672_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11376_ _05304_ net458 _05629_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10327_ _05040_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13115_ clknet_leaf_131_clk _00573_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ clknet_leaf_23_clk _00504_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[19\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10258_ _05002_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10189_ _04877_ net421 _04952_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06420_ _01337_ rvsingle.dp.rf.rf\[22\]\[29\] _01302_ VGND VGND VPWR VPWR _01342_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06351_ rvsingle.dp.rf.rf\[16\]\[29\] rvsingle.dp.rf.rf\[17\]\[29\] rvsingle.dp.rf.rf\[18\]\[29\]
+ rvsingle.dp.rf.rf\[19\]\[29\] _01139_ _01261_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09070_ _01330_ rvsingle.dp.rf.rf\[6\]\[26\] VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06282_ rvsingle.dp.rf.rf\[8\]\[30\] rvsingle.dp.rf.rf\[9\]\[30\] rvsingle.dp.rf.rf\[10\]\[30\]
+ rvsingle.dp.rf.rf\[11\]\[30\] _01196_ _01203_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08021_ _02440_ rvsingle.dp.rf.rf\[10\]\[0\] _01243_ VGND VGND VPWR VPWR _02942_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold702 rvsingle.dp.rf.rf\[16\]\[3\] VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 rvsingle.dp.rf.rf\[13\]\[18\] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold724 rvsingle.dp.rf.rf\[15\]\[7\] VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold735 rvsingle.dp.rf.rf\[22\]\[1\] VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold746 rvsingle.dp.rf.rf\[18\]\[26\] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold757 rvsingle.dp.rf.rf\[29\]\[6\] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 rvsingle.dp.rf.rf\[9\]\[6\] VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold779 rvsingle.dp.rf.rf\[23\]\[6\] VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09972_ DataAdr[11] ReadData[11] _04750_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08923_ _01138_ rvsingle.dp.rf.rf\[20\]\[25\] VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08854_ _02266_ _03759_ _03774_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__o21bai_4
X_07805_ _01520_ _02722_ _02723_ _01111_ _02725_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__o311ai_2
X_08785_ rvsingle.dp.rf.rf\[20\]\[15\] rvsingle.dp.rf.rf\[21\]\[15\] rvsingle.dp.rf.rf\[22\]\[15\]
+ rvsingle.dp.rf.rf\[23\]\[15\] _01691_ _01244_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__mux4_2
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ _02644_ _02656_ _01145_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__nand3_2
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07667_ _01349_ rvsingle.dp.rf.rf\[10\]\[5\] VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09406_ _03561_ _01185_ _02261_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06618_ _01086_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__buf_6
X_07598_ rvsingle.dp.rf.rf\[29\]\[4\] _01267_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09337_ _02184_ _04250_ _04251_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__nand3b_2
X_06549_ _01454_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09268_ _01250_ _04061_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08219_ _01201_ _01351_ _03124_ _03139_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09199_ _01250_ _04063_ _04116_ _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_105_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11230_ _05554_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11161_ _05516_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__clkbuf_1
X_10112_ _04907_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__clkbuf_2
X_11092_ _05479_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__clkbuf_1
X_10043_ _04848_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__clkbuf_1
Xhold40 rvsingle.dp.rf.rf\[22\]\[31\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 rvsingle.dp.rf.rf\[19\]\[31\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 rvsingle.dp.rf.rf\[3\]\[31\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 rvsingle.dp.rf.rf\[1\]\[31\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 rvsingle.dp.rf.rf\[26\]\[31\] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 rvsingle.dp.rf.rf\[7\]\[14\] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11994_ _05757_ rvsingle.dp.rf.rf\[4\]\[23\] _05960_ VGND VGND VPWR VPWR _05964_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10945_ _05399_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10876_ _04877_ net296 _05319_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12615_ clknet_leaf_104_clk _00073_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[22\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12546_ clknet_leaf_126_clk _01030_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12477_ clknet_leaf_146_clk _00961_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[26\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_4 DataAdr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11428_ _05291_ net723 _05657_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11359_ _05476_ net785 _05618_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ clknet_leaf_111_clk _00487_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[11\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08570_ _01469_ rvsingle.dp.rf.rf\[8\]\[12\] VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07521_ _01707_ rvsingle.dp.rf.rf\[4\]\[6\] VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07452_ _01065_ _02318_ _01870_ _02319_ _02372_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_146_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06403_ rvsingle.dp.rf.rf\[24\]\[29\] rvsingle.dp.rf.rf\[25\]\[29\] rvsingle.dp.rf.rf\[26\]\[29\]
+ rvsingle.dp.rf.rf\[27\]\[29\] _01194_ _01303_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07383_ _01468_ rvsingle.dp.rf.rf\[18\]\[7\] VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09122_ rvsingle.dp.rf.rf\[28\]\[26\] rvsingle.dp.rf.rf\[29\]\[26\] rvsingle.dp.rf.rf\[30\]\[26\]
+ rvsingle.dp.rf.rf\[31\]\[26\] _01643_ _01491_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__mux4_1
X_06334_ _01256_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__buf_4
XFILLER_0_161_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09053_ _01744_ rvsingle.dp.rf.rf\[14\]\[27\] _01648_ VGND VGND VPWR VPWR _03973_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06265_ _01187_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_142_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08004_ _02921_ _02922_ _01172_ _02924_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold510 rvsingle.dp.rf.rf\[18\]\[25\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06196_ _01107_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__clkbuf_4
Xhold521 rvsingle.dp.rf.rf\[21\]\[18\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold532 rvsingle.dp.rf.rf\[0\]\[15\] VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 rvsingle.dp.rf.rf\[6\]\[17\] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 rvsingle.dp.rf.rf\[0\]\[13\] VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 rvsingle.dp.rf.rf\[27\]\[16\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold576 rvsingle.dp.rf.rf\[4\]\[11\] VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 rvsingle.dp.rf.rf\[10\]\[22\] VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 rvsingle.dp.rf.rf\[10\]\[4\] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _04774_ net406 _04741_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__mux2_1
X_08906_ _03803_ _03825_ _03826_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__nand3b_2
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _01078_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__buf_4
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _03745_ _03754_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__o21ai_2
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _03685_ _03686_ _02351_ _03688_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__o211ai_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ rvsingle.dp.rf.rf\[25\]\[5\] _01877_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__and2b_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _03608_ _03619_ _01146_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__nand3_4
XFILLER_0_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10730_ _04909_ _04913_ _05232_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10661_ _04918_ _04922_ _05057_ _04916_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__and4b_2
XFILLER_0_94_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12400_ clknet_leaf_53_clk _00884_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[28\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13380_ clknet_leaf_91_clk _00808_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[5\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_994 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10592_ _05193_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__buf_6
XFILLER_0_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12331_ _04823_ net373 _06110_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12262_ _05474_ _05847_ _06077_ net82 VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_105_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11213_ _05545_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__clkbuf_1
X_12193_ _06062_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
X_11144_ _05507_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11075_ _05209_ net692 _05469_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10026_ _04833_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11977_ _05955_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10928_ _05209_ net817 _05387_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10859_ _05347_ _05069_ _05068_ _05320_ net12 VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12529_ clknet_leaf_49_clk _01013_ VGND VGND VPWR VPWR rvsingle.dp.rf.rf\[24\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06952_ _01862_ rvsingle.dp.rf.rf\[28\]\[22\] VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__or2_1
X_09740_ _04578_ _04579_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__xor2_1
.ends

